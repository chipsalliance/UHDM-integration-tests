module bsg_nor3(a_i, b_i, c_i, o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  input [15:0] a_i;
  wire [15:0] a_i;
  input [15:0] b_i;
  wire [15:0] b_i;
  input [15:0] c_i;
  wire [15:0] c_i;
  output [15:0] o;
  wire [15:0] o;
  assign _00_ = ~(b_i[0] | a_i[0]);
  assign o[0] = _00_ & ~(c_i[0]);
  assign _01_ = ~(b_i[1] | a_i[1]);
  assign o[1] = _01_ & ~(c_i[1]);
  assign _02_ = ~(b_i[2] | a_i[2]);
  assign o[2] = _02_ & ~(c_i[2]);
  assign _03_ = ~(b_i[3] | a_i[3]);
  assign o[3] = _03_ & ~(c_i[3]);
  assign _04_ = ~(b_i[4] | a_i[4]);
  assign o[4] = _04_ & ~(c_i[4]);
  assign _05_ = ~(b_i[5] | a_i[5]);
  assign o[5] = _05_ & ~(c_i[5]);
  assign _06_ = ~(b_i[6] | a_i[6]);
  assign o[6] = _06_ & ~(c_i[6]);
  assign _07_ = ~(b_i[7] | a_i[7]);
  assign o[7] = _07_ & ~(c_i[7]);
  assign _08_ = ~(b_i[8] | a_i[8]);
  assign o[8] = _08_ & ~(c_i[8]);
  assign _09_ = ~(b_i[9] | a_i[9]);
  assign o[9] = _09_ & ~(c_i[9]);
  assign _10_ = ~(b_i[10] | a_i[10]);
  assign o[10] = _10_ & ~(c_i[10]);
  assign _11_ = ~(b_i[11] | a_i[11]);
  assign o[11] = _11_ & ~(c_i[11]);
  assign _12_ = ~(b_i[12] | a_i[12]);
  assign o[12] = _12_ & ~(c_i[12]);
  assign _13_ = ~(b_i[13] | a_i[13]);
  assign o[13] = _13_ & ~(c_i[13]);
  assign _14_ = ~(b_i[14] | a_i[14]);
  assign o[14] = _14_ & ~(c_i[14]);
  assign _15_ = ~(b_i[15] | a_i[15]);
  assign o[15] = _15_ & ~(c_i[15]);
endmodule
