module bsg_clkbuf(i, o);
  input [15:0] i;
  wire [15:0] i;
  output [15:0] o;
  wire [15:0] o;
  assign o = i;
endmodule
