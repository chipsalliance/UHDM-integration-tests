module bsg_compare_and_swap(data_i, swap_on_equal_i, data_o, swapped_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  input [31:0] data_i;
  wire [31:0] data_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire gt;
  input swap_on_equal_i;
  wire swap_on_equal_i;
  output swapped_o;
  wire swapped_o;
  assign _043_ = data_i[15] & ~(data_i[31]);
  assign _044_ = ~(data_i[15] ^ data_i[31]);
  assign _045_ = data_i[30] | ~(data_i[14]);
  assign _046_ = _044_ & ~(_045_);
  assign _047_ = _046_ | _043_;
  assign _048_ = data_i[14] ^ data_i[30];
  assign _049_ = _044_ & ~(_048_);
  assign _050_ = data_i[29] | ~(data_i[13]);
  assign _051_ = data_i[13] ^ data_i[29];
  assign _052_ = data_i[12] & ~(data_i[28]);
  assign _053_ = _052_ & ~(_051_);
  assign _054_ = _050_ & ~(_053_);
  assign _055_ = _049_ & ~(_054_);
  assign _056_ = _055_ | _047_;
  assign _057_ = data_i[12] ^ data_i[28];
  assign _058_ = _057_ | _051_;
  assign _059_ = _049_ & ~(_058_);
  assign _060_ = data_i[27] | ~(data_i[11]);
  assign _061_ = ~(data_i[11] ^ data_i[27]);
  assign _062_ = data_i[26] | ~(data_i[10]);
  assign _063_ = _061_ & ~(_062_);
  assign _064_ = _060_ & ~(_063_);
  assign _065_ = data_i[10] ^ data_i[26];
  assign _066_ = _065_ | ~(_061_);
  assign _067_ = data_i[25] | ~(data_i[9]);
  assign _068_ = data_i[9] ^ data_i[25];
  assign _069_ = data_i[8] & ~(data_i[24]);
  assign _070_ = _069_ & ~(_068_);
  assign _071_ = _070_ | ~(_067_);
  assign _072_ = _071_ & ~(_066_);
  assign _073_ = _064_ & ~(_072_);
  assign _074_ = _059_ & ~(_073_);
  assign _075_ = _074_ | _056_;
  assign _076_ = data_i[8] ^ data_i[24];
  assign _000_ = _076_ | _068_;
  assign _001_ = _000_ | _066_;
  assign _002_ = _059_ & ~(_001_);
  assign _003_ = data_i[23] | ~(data_i[7]);
  assign _004_ = ~(data_i[7] ^ data_i[23]);
  assign _005_ = data_i[22] | ~(data_i[6]);
  assign _006_ = _004_ & ~(_005_);
  assign _007_ = _003_ & ~(_006_);
  assign _008_ = data_i[6] ^ data_i[22];
  assign _009_ = _004_ & ~(_008_);
  assign _010_ = data_i[21] | ~(data_i[5]);
  assign _011_ = data_i[5] ^ data_i[21];
  assign _012_ = data_i[4] & ~(data_i[20]);
  assign _013_ = _012_ & ~(_011_);
  assign _014_ = _010_ & ~(_013_);
  assign _015_ = _009_ & ~(_014_);
  assign _016_ = _007_ & ~(_015_);
  assign _017_ = data_i[4] ^ data_i[20];
  assign _018_ = _017_ | _011_;
  assign _019_ = _018_ | ~(_009_);
  assign _020_ = data_i[19] | ~(data_i[3]);
  assign _021_ = ~(data_i[3] ^ data_i[19]);
  assign _022_ = data_i[18] | ~(data_i[2]);
  assign _023_ = _021_ & ~(_022_);
  assign _024_ = _020_ & ~(_023_);
  assign _025_ = data_i[2] ^ data_i[18];
  assign _026_ = _025_ | ~(_021_);
  assign _027_ = data_i[17] | ~(data_i[1]);
  assign _028_ = data_i[1] ^ data_i[17];
  assign _029_ = data_i[0] | ~(data_i[16]);
  assign _030_ = _029_ & ~(_028_);
  assign _031_ = _030_ | ~(_027_);
  assign _032_ = _031_ & ~(_026_);
  assign _033_ = _032_ | ~(_024_);
  assign _034_ = _033_ & ~(_019_);
  assign _035_ = _016_ & ~(_034_);
  assign _036_ = _002_ & ~(_035_);
  assign _037_ = _036_ | _075_;
  assign _038_ = data_i[0] ^ data_i[16];
  assign _039_ = _038_ | _028_;
  assign _040_ = _039_ | _026_;
  assign _041_ = _040_ | _019_;
  assign _042_ = _002_ & ~(_041_);
  assign swapped_o = _037_ & ~(_042_);
  assign data_o[0] = swapped_o ? data_i[16] : data_i[0];
  assign data_o[1] = swapped_o ? data_i[17] : data_i[1];
  assign data_o[2] = swapped_o ? data_i[18] : data_i[2];
  assign data_o[3] = swapped_o ? data_i[19] : data_i[3];
  assign data_o[4] = swapped_o ? data_i[20] : data_i[4];
  assign data_o[5] = swapped_o ? data_i[21] : data_i[5];
  assign data_o[6] = swapped_o ? data_i[22] : data_i[6];
  assign data_o[7] = swapped_o ? data_i[23] : data_i[7];
  assign data_o[8] = swapped_o ? data_i[24] : data_i[8];
  assign data_o[9] = swapped_o ? data_i[25] : data_i[9];
  assign data_o[10] = swapped_o ? data_i[26] : data_i[10];
  assign data_o[11] = swapped_o ? data_i[27] : data_i[11];
  assign data_o[12] = swapped_o ? data_i[28] : data_i[12];
  assign data_o[13] = swapped_o ? data_i[29] : data_i[13];
  assign data_o[14] = swapped_o ? data_i[30] : data_i[14];
  assign data_o[15] = swapped_o ? data_i[31] : data_i[15];
  assign data_o[16] = swapped_o ? data_i[0] : data_i[16];
  assign data_o[17] = swapped_o ? data_i[1] : data_i[17];
  assign data_o[18] = swapped_o ? data_i[2] : data_i[18];
  assign data_o[19] = swapped_o ? data_i[3] : data_i[19];
  assign data_o[20] = swapped_o ? data_i[4] : data_i[20];
  assign data_o[21] = swapped_o ? data_i[5] : data_i[21];
  assign data_o[22] = swapped_o ? data_i[6] : data_i[22];
  assign data_o[23] = swapped_o ? data_i[7] : data_i[23];
  assign data_o[24] = swapped_o ? data_i[8] : data_i[24];
  assign data_o[25] = swapped_o ? data_i[9] : data_i[25];
  assign data_o[26] = swapped_o ? data_i[10] : data_i[26];
  assign data_o[27] = swapped_o ? data_i[11] : data_i[27];
  assign data_o[28] = swapped_o ? data_i[12] : data_i[28];
  assign data_o[29] = swapped_o ? data_i[13] : data_i[29];
  assign data_o[30] = swapped_o ? data_i[14] : data_i[30];
  assign data_o[31] = swapped_o ? data_i[15] : data_i[31];
  assign gt = swapped_o;
endmodule
