module bsg_swap(data_i, swap_i, data_o);
  input [31:0] data_i;
  wire [31:0] data_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  input swap_i;
  wire swap_i;
  assign data_o[21] = swap_i ? data_i[5] : data_i[21];
  assign data_o[22] = swap_i ? data_i[6] : data_i[22];
  assign data_o[23] = swap_i ? data_i[7] : data_i[23];
  assign data_o[24] = swap_i ? data_i[8] : data_i[24];
  assign data_o[25] = swap_i ? data_i[9] : data_i[25];
  assign data_o[26] = swap_i ? data_i[10] : data_i[26];
  assign data_o[27] = swap_i ? data_i[11] : data_i[27];
  assign data_o[28] = swap_i ? data_i[12] : data_i[28];
  assign data_o[29] = swap_i ? data_i[13] : data_i[29];
  assign data_o[30] = swap_i ? data_i[14] : data_i[30];
  assign data_o[31] = swap_i ? data_i[15] : data_i[31];
  assign data_o[0] = swap_i ? data_i[16] : data_i[0];
  assign data_o[1] = swap_i ? data_i[17] : data_i[1];
  assign data_o[2] = swap_i ? data_i[18] : data_i[2];
  assign data_o[3] = swap_i ? data_i[19] : data_i[3];
  assign data_o[4] = swap_i ? data_i[20] : data_i[4];
  assign data_o[5] = swap_i ? data_i[21] : data_i[5];
  assign data_o[6] = swap_i ? data_i[22] : data_i[6];
  assign data_o[7] = swap_i ? data_i[23] : data_i[7];
  assign data_o[8] = swap_i ? data_i[24] : data_i[8];
  assign data_o[9] = swap_i ? data_i[25] : data_i[9];
  assign data_o[10] = swap_i ? data_i[26] : data_i[10];
  assign data_o[11] = swap_i ? data_i[27] : data_i[11];
  assign data_o[12] = swap_i ? data_i[28] : data_i[12];
  assign data_o[13] = swap_i ? data_i[29] : data_i[13];
  assign data_o[14] = swap_i ? data_i[30] : data_i[14];
  assign data_o[15] = swap_i ? data_i[31] : data_i[15];
  assign data_o[16] = swap_i ? data_i[0] : data_i[16];
  assign data_o[17] = swap_i ? data_i[1] : data_i[17];
  assign data_o[18] = swap_i ? data_i[2] : data_i[18];
  assign data_o[19] = swap_i ? data_i[3] : data_i[19];
  assign data_o[20] = swap_i ? data_i[4] : data_i[20];
endmodule
