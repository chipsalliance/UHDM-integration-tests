module bsg_priority_encode_one_hot_out(i, o, v_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  input [15:0] i;
  wire [15:0] i;
  wire [15:0] \nw1.scan.i ;
  wire [15:0] \nw1.scan.o ;
  wire [15:0] \nw1.scan.scanN.row[0].fill ;
  wire [15:0] \nw1.scan.scanN.row[0].shifted ;
  wire [15:0] \nw1.scan.scanN.row[1].fill ;
  wire [15:0] \nw1.scan.scanN.row[1].shifted ;
  wire [15:0] \nw1.scan.scanN.row[2].fill ;
  wire [15:0] \nw1.scan.scanN.row[2].shifted ;
  wire [15:0] \nw1.scan.scanN.row[3].fill ;
  wire [15:0] \nw1.scan.scanN.row[3].shifted ;
  wire [79:0] \nw1.scan.t ;
  output [15:0] o;
  wire [15:0] o;
  wire [15:0] scan_lo;
  output v_o;
  wire v_o;
  assign _000_ = i[1] | i[0];
  assign _001_ = i[3] | i[2];
  assign _002_ = _001_ | _000_;
  assign _003_ = i[5] | i[4];
  assign _004_ = i[7] | i[6];
  assign _005_ = _004_ | _003_;
  assign _006_ = _005_ | _002_;
  assign _007_ = i[9] | i[8];
  assign _008_ = i[11] | i[10];
  assign _009_ = _008_ | _007_;
  assign _010_ = i[13] | i[12];
  assign _011_ = i[14] | i[15];
  assign _012_ = _011_ | _010_;
  assign _013_ = _012_ | _009_;
  assign v_o = _013_ | _006_;
  assign _014_ = i[2] | i[1];
  assign _015_ = i[4] | i[3];
  assign _016_ = _015_ | _014_;
  assign _017_ = i[6] | i[5];
  assign _018_ = i[8] | i[7];
  assign _019_ = _018_ | _017_;
  assign _020_ = _019_ | _016_;
  assign _021_ = i[10] | i[9];
  assign _022_ = i[12] | i[11];
  assign _023_ = _022_ | _021_;
  assign _024_ = i[14] | i[13];
  assign _025_ = _024_ | i[15];
  assign _026_ = _025_ | _023_;
  assign _027_ = _026_ | _020_;
  assign o[0] = v_o & ~(_027_);
  assign _028_ = _003_ | _001_;
  assign _029_ = _007_ | _004_;
  assign _030_ = _029_ | _028_;
  assign _031_ = _010_ | _008_;
  assign _032_ = _031_ | _011_;
  assign _033_ = _032_ | _030_;
  assign o[1] = _027_ & ~(_033_);
  assign _034_ = _017_ | _015_;
  assign _035_ = _021_ | _018_;
  assign _036_ = _035_ | _034_;
  assign _037_ = _024_ | _022_;
  assign _038_ = _037_ | i[15];
  assign _039_ = _038_ | _036_;
  assign o[2] = _033_ & ~(_039_);
  assign _040_ = _009_ | _005_;
  assign _041_ = _040_ | _012_;
  assign o[3] = _039_ & ~(_041_);
  assign _042_ = _023_ | _019_;
  assign _043_ = _042_ | _025_;
  assign o[4] = _041_ & ~(_043_);
  assign _044_ = _031_ | _029_;
  assign _045_ = _044_ | _011_;
  assign o[5] = _043_ & ~(_045_);
  assign _046_ = _037_ | _035_;
  assign _047_ = _046_ | i[15];
  assign o[6] = _045_ & ~(_047_);
  assign o[7] = _047_ & ~(_013_);
  assign o[8] = _013_ & ~(_026_);
  assign o[9] = _026_ & ~(_032_);
  assign o[10] = _032_ & ~(_038_);
  assign o[11] = _038_ & ~(_012_);
  assign o[12] = _012_ & ~(_025_);
  assign o[13] = _025_ & ~(_011_);
  assign o[14] = i[14] & ~(i[15]);
  assign \nw1.scan.i  = i;
  assign { \nw1.scan.o [15], \nw1.scan.o [0] } = { i[15], v_o };
  assign \nw1.scan.scanN.row[0].fill  = 16'h0000;
  assign \nw1.scan.scanN.row[0].shifted  = { 1'h0, i[15:1] };
  assign \nw1.scan.scanN.row[1].fill  = 16'h0000;
  assign \nw1.scan.scanN.row[1].shifted [15:12] = { 2'h0, i[15], \nw1.scan.o [14] };
  assign \nw1.scan.scanN.row[2].fill  = 16'h0000;
  assign \nw1.scan.scanN.row[2].shifted [15:8] = { 4'h0, i[15], \nw1.scan.o [14:12] };
  assign \nw1.scan.scanN.row[3].fill  = 16'h0000;
  assign \nw1.scan.scanN.row[3].shifted  = { 8'h00, i[15], \nw1.scan.o [14:8] };
  assign { \nw1.scan.t [79:56], \nw1.scan.t [47:36], \nw1.scan.t [31:18], \nw1.scan.t [15:0] } = { i[15], \nw1.scan.o [14:1], v_o, i[15], \nw1.scan.o [14:8], i[15], \nw1.scan.o [14:12], \nw1.scan.scanN.row[2].shifted [7:0], i[15], \nw1.scan.o [14], \nw1.scan.scanN.row[1].shifted [11:0], i };
  assign o[15] = i[15];
  assign scan_lo = { i[15], \nw1.scan.o [14:1], v_o };
endmodule
