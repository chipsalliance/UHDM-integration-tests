module top;
  import flash_ctrl_pkg::*;
endmodule
