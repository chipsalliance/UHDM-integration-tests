module bsg_fsb_murn_gateway(clk_i, reset_i, v_i, data_i, ready_o, v_o, ready_i, node_en_r_o, node_reset_r_o);
  input clk_i;
  wire clk_i;
  input [15:0] data_i;
  wire [15:0] data_i;
  wire [21:0] \genblk1.data_RPT ;
  wire \genblk1.for_switch ;
  wire \genblk1.for_this_node ;
  wire \genblk1.id_match ;
  wire \genblk1.node_en_n ;
  wire \genblk1.node_en_r ;
  wire \genblk1.node_reset_n ;
  wire \genblk1.node_reset_r ;
  output node_en_r_o;
  wire node_en_r_o;
  output node_reset_r_o;
  wire node_reset_r_o;
  input ready_i;
  wire ready_i;
  output ready_o;
  wire ready_o;
  input reset_i;
  wire reset_i;
  input v_i;
  wire v_i;
  output v_o;
  wire v_o;
  assign \genblk1.data_RPT  = { 6'h00, data_i };
  assign \genblk1.for_switch  = 1'h0;
  assign \genblk1.for_this_node  = 1'h0;
  assign \genblk1.id_match  = 1'h0;
  assign \genblk1.node_en_n  = 1'h0;
  assign \genblk1.node_en_r  = 1'h0;
  assign \genblk1.node_reset_n  = 1'h1;
  assign \genblk1.node_reset_r  = 1'h1;
  assign node_en_r_o = 1'h0;
  assign node_reset_r_o = 1'h1;
  assign ready_o = v_i;
  assign v_o = 1'h0;
endmodule
