module bsg_priority_encode(i, addr_o, v_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire [15:0] \a.i ;
  wire [15:0] \a.nw1.scan.i ;
  wire [15:0] \a.nw1.scan.o ;
  wire [15:0] \a.nw1.scan.scanN.row[0].fill ;
  wire [15:0] \a.nw1.scan.scanN.row[0].shifted ;
  wire [15:0] \a.nw1.scan.scanN.row[1].fill ;
  wire [15:0] \a.nw1.scan.scanN.row[1].shifted ;
  wire [15:0] \a.nw1.scan.scanN.row[2].fill ;
  wire [15:0] \a.nw1.scan.scanN.row[2].shifted ;
  wire [15:0] \a.nw1.scan.scanN.row[3].fill ;
  wire [15:0] \a.nw1.scan.scanN.row[3].shifted ;
  wire [79:0] \a.nw1.scan.t ;
  wire [15:0] \a.o ;
  wire [15:0] \a.scan_lo ;
  wire \a.v_o ;
  output [3:0] addr_o;
  wire [3:0] addr_o;
  wire [79:0] \b.addr ;
  wire [3:0] \b.addr_o ;
  wire [15:0] \b.i ;
  wire [1:0] \b.rof[1].rof1[0].vs ;
  wire [1:0] \b.rof[1].rof1[1].vs ;
  wire [1:0] \b.rof[1].rof1[2].vs ;
  wire [1:0] \b.rof[1].rof1[3].vs ;
  wire [1:0] \b.rof[1].rof1[4].vs ;
  wire [1:0] \b.rof[1].rof1[5].vs ;
  wire [1:0] \b.rof[1].rof1[6].vs ;
  wire [1:0] \b.rof[1].rof1[7].vs ;
  wire [1:0] \b.rof[2].rof1[0].vs ;
  wire [1:0] \b.rof[2].rof1[1].vs ;
  wire [1:0] \b.rof[2].rof1[2].vs ;
  wire [1:0] \b.rof[2].rof1[3].vs ;
  wire [1:0] \b.rof[3].rof1[0].vs ;
  wire [1:0] \b.rof[3].rof1[1].vs ;
  wire [1:0] \b.rof[4].rof1[0].vs ;
  wire [79:0] \b.v ;
  wire \b.v_o ;
  wire [14:0] enc_lo;
  input [15:0] i;
  wire [15:0] i;
  output v_o;
  wire v_o;
  assign _002_ = i[1] | i[0];
  assign _003_ = i[3] | i[2];
  assign _004_ = _003_ | _002_;
  assign _005_ = i[5] | i[4];
  assign _006_ = i[7] | i[6];
  assign _007_ = _006_ | _005_;
  assign _008_ = _007_ | _004_;
  assign _009_ = i[9] | i[8];
  assign _010_ = i[11] | i[10];
  assign _011_ = _010_ | _009_;
  assign _012_ = i[13] | i[12];
  assign _013_ = i[14] | i[15];
  assign _014_ = _013_ | _012_;
  assign _015_ = _014_ | _011_;
  assign v_o = _015_ | _008_;
  assign _016_ = ~(i[2] | i[1]);
  assign _017_ = i[4] | i[3];
  assign _018_ = _016_ & ~(_017_);
  assign _019_ = i[6] | i[5];
  assign _020_ = i[8] | i[7];
  assign _021_ = _020_ | _019_;
  assign _022_ = _018_ & ~(_021_);
  assign _023_ = i[10] | i[9];
  assign _024_ = i[12] | i[11];
  assign _025_ = _024_ | _023_;
  assign _026_ = i[14] | i[13];
  assign _027_ = _026_ | i[15];
  assign _028_ = _027_ | _025_;
  assign _029_ = _022_ & ~(_028_);
  assign _030_ = ~(_005_ | _003_);
  assign _031_ = _009_ | _006_;
  assign _032_ = _030_ & ~(_031_);
  assign _033_ = _012_ | _010_;
  assign _034_ = _033_ | _013_;
  assign _035_ = _032_ & ~(_034_);
  assign _036_ = _029_ ? v_o : _035_;
  assign _037_ = ~(_019_ | _017_);
  assign _038_ = _023_ | _020_;
  assign _039_ = _037_ & ~(_038_);
  assign _040_ = _026_ | _024_;
  assign _041_ = _040_ | i[15];
  assign _042_ = _039_ & ~(_041_);
  assign _043_ = _011_ | _007_;
  assign _044_ = _043_ | _014_;
  assign _045_ = _042_ ? _035_ : _044_;
  assign _046_ = _036_ | ~(_045_);
  assign _047_ = _025_ | _021_;
  assign _048_ = ~(_047_ | _027_);
  assign _049_ = _033_ | _031_;
  assign _050_ = ~(_049_ | _013_);
  assign _051_ = _048_ ? _044_ : _050_;
  assign _052_ = _040_ | _038_;
  assign _053_ = _052_ | i[15];
  assign _054_ = _053_ ? _015_ : _050_;
  assign _055_ = _051_ | ~(_054_);
  assign addr_o[3] = _055_ | _046_;
  assign _056_ = _029_ & v_o;
  assign _057_ = _042_ & ~(_035_);
  assign _058_ = _057_ | _056_;
  assign _059_ = _048_ & _044_;
  assign _060_ = ~(_053_ | _050_);
  assign _061_ = _060_ | _059_;
  assign _062_ = _061_ | _058_;
  assign _063_ = _015_ & ~(_028_);
  assign _064_ = _034_ & ~(_041_);
  assign _065_ = _064_ | _063_;
  assign _066_ = _014_ & ~(_027_);
  assign _067_ = i[14] & ~(i[15]);
  assign _068_ = _067_ | _066_;
  assign _069_ = _068_ | _065_;
  assign addr_o[0] = _069_ | _062_;
  assign _070_ = _051_ | _036_;
  assign _071_ = ~_034_;
  assign _072_ = _028_ ? _071_ : _015_;
  assign _073_ = ~_013_;
  assign _074_ = _027_ ? _073_ : _014_;
  assign _075_ = _074_ | _072_;
  assign addr_o[1] = _075_ | _070_;
  assign _000_ = _041_ ? _014_ : _071_;
  assign _001_ = _072_ | ~(_000_);
  assign addr_o[2] = _001_ | _046_;
  assign \a.i  = i;
  assign \a.nw1.scan.i  = i;
  assign { \a.nw1.scan.o [15], \a.nw1.scan.o [0] } = { i[15], v_o };
  assign \a.nw1.scan.scanN.row[0].fill  = 16'h0000;
  assign \a.nw1.scan.scanN.row[0].shifted  = { 1'h0, i[15:1] };
  assign \a.nw1.scan.scanN.row[1].fill  = 16'h0000;
  assign \a.nw1.scan.scanN.row[1].shifted [15:12] = { 2'h0, i[15], \a.nw1.scan.o [14] };
  assign \a.nw1.scan.scanN.row[2].fill  = 16'h0000;
  assign \a.nw1.scan.scanN.row[2].shifted [15:8] = { 4'h0, i[15], \a.nw1.scan.o [14:12] };
  assign \a.nw1.scan.scanN.row[3].fill  = 16'h0000;
  assign \a.nw1.scan.scanN.row[3].shifted  = { 8'h00, i[15], \a.nw1.scan.o [14:8] };
  assign { \a.nw1.scan.t [79:56], \a.nw1.scan.t [47:36], \a.nw1.scan.t [31:18], \a.nw1.scan.t [15:0] } = { i[15], \a.nw1.scan.o [14:1], v_o, i[15], \a.nw1.scan.o [14:8], i[15], \a.nw1.scan.o [14:12], \a.nw1.scan.scanN.row[2].shifted [7:0], i[15], \a.nw1.scan.o [14], \a.nw1.scan.scanN.row[1].shifted [11:0], i };
  assign \a.o [15] = 1'hx;
  assign \a.scan_lo  = { i[15], \a.nw1.scan.o [14:1], v_o };
  assign \a.v_o  = v_o;
  assign { \b.addr [79:59], \b.addr [55:51], \b.addr [47:46], \b.addr [43:42], \b.addr [39:38], \b.addr [35:34], \b.addr [31:0] } = { 12'hxxx, addr_o, 19'hxxxxx, \a.o [14], 1'hx, \a.o [12], 1'hx, \a.o [10], 1'hx, \a.o [8], 1'hx, \a.o [6], 1'hx, \a.o [4], 1'hx, \a.o [2], 1'hx, \a.o [0], 16'h0000 };
  assign \b.addr_o  = addr_o;
  assign \b.i  = { 1'hx, \a.o [14:0] };
  assign \b.rof[1].rof1[0].vs  = \a.o [1:0];
  assign \b.rof[1].rof1[1].vs  = \a.o [3:2];
  assign \b.rof[1].rof1[2].vs  = \a.o [5:4];
  assign \b.rof[1].rof1[3].vs  = \a.o [7:6];
  assign \b.rof[1].rof1[4].vs  = \a.o [9:8];
  assign \b.rof[1].rof1[5].vs  = \a.o [11:10];
  assign \b.rof[1].rof1[6].vs  = \a.o [13:12];
  assign \b.rof[1].rof1[7].vs  = { 1'hx, \a.o [14] };
  assign \b.rof[2].rof1[0].vs  = { 1'hx, \b.addr [33] };
  assign \b.rof[2].rof1[1].vs  = { 1'hx, \b.addr [37] };
  assign \b.rof[2].rof1[2].vs  = { 1'hx, \b.addr [41] };
  assign \b.rof[2].rof1[3].vs  = { 1'hx, \b.addr [45] };
  assign \b.rof[3].rof1[0].vs  = { 1'hx, \b.addr [50] };
  assign \b.rof[3].rof1[1].vs  = { 1'hx, \b.addr [58] };
  assign \b.rof[4].rof1[0].vs  = { 1'hx, addr_o[3] };
  assign \b.v  = { 31'hxxxxxxxx, addr_o[3], 7'hxx, \b.addr [58], 7'hxx, \b.addr [50], 3'hx, \b.addr [45], 3'hx, \b.addr [41], 3'hx, \b.addr [37], 3'hx, \b.addr [33], 1'hx, \a.o [14:0] };
  assign \b.v_o  = 1'hx;
  assign enc_lo = \a.o [14:0];
endmodule
