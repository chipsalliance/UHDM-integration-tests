module bsg_tielo(o);
  output [15:0] o;
  wire [15:0] o;
  assign o = 16'h0000;
endmodule
