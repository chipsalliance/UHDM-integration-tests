module top(output logic o);
   assign o = logic'(1);
endmodule
