module bsg_lru_pseudo_tree_decode(way_id_i, data_o, mask_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  output [14:0] data_o;
  wire [14:0] data_o;
  output [14:0] mask_o;
  wire [14:0] mask_o;
  input [3:0] way_id_i;
  wire [3:0] way_id_i;
  assign data_o[0] = ~way_id_i[3];
  assign _00_ = way_id_i[2] | way_id_i[3];
  assign data_o[1] = ~_00_;
  assign _01_ = way_id_i[2] | ~(way_id_i[3]);
  assign data_o[2] = ~_01_;
  assign _02_ = way_id_i[3] | ~(way_id_i[2]);
  assign mask_o[4] = ~_02_;
  assign _03_ = ~(way_id_i[2] & way_id_i[3]);
  assign mask_o[6] = ~_03_;
  assign _04_ = ~way_id_i[1];
  assign data_o[3] = _04_ & ~(_00_);
  assign data_o[7] = data_o[3] & ~(way_id_i[0]);
  assign mask_o[8] = way_id_i[1] & ~(_00_);
  assign data_o[8] = mask_o[8] & ~(way_id_i[0]);
  assign data_o[4] = _04_ & ~(_02_);
  assign data_o[9] = data_o[4] & ~(way_id_i[0]);
  assign mask_o[10] = way_id_i[1] & ~(_02_);
  assign data_o[10] = mask_o[10] & ~(way_id_i[0]);
  assign data_o[5] = _04_ & ~(_01_);
  assign data_o[11] = data_o[5] & ~(way_id_i[0]);
  assign mask_o[12] = way_id_i[1] & ~(_01_);
  assign data_o[12] = mask_o[12] & ~(way_id_i[0]);
  assign data_o[6] = _04_ & ~(_03_);
  assign data_o[13] = data_o[6] & ~(way_id_i[0]);
  assign mask_o[14] = way_id_i[1] & ~(_03_);
  assign data_o[14] = mask_o[14] & ~(way_id_i[0]);
  assign { mask_o[13], mask_o[11], mask_o[9], mask_o[7], mask_o[5], mask_o[3:0] } = { data_o[6:1], way_id_i[3], data_o[0], 1'h1 };
endmodule
