module bsg_round_robin_2_to_2(clk_i, reset_i, data_i, v_i, ready_o, data_o, v_o, ready_i);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  input clk_i;
  wire clk_i;
  input [31:0] data_i;
  wire [31:0] data_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  reg head_r;
  input [1:0] ready_i;
  wire [1:0] ready_i;
  output [1:0] ready_o;
  wire [1:0] ready_o;
  input reset_i;
  wire reset_i;
  input [1:0] v_i;
  wire [1:0] v_i;
  output [1:0] v_o;
  wire [1:0] v_o;
  assign ready_o[0] = head_r ? ready_i[1] : ready_i[0];
  assign _00_ = ~(ready_o[0] & v_i[0]);
  assign ready_o[1] = head_r ? ready_i[0] : ready_i[1];
  assign _01_ = ready_o[1] & v_i[1];
  assign _02_ = ~(_01_ ^ _00_);
  assign _03_ = _02_ ^ head_r;
  assign data_o[11] = head_r ? data_i[27] : data_i[11];
  assign data_o[12] = head_r ? data_i[28] : data_i[12];
  assign data_o[13] = head_r ? data_i[29] : data_i[13];
  assign data_o[14] = head_r ? data_i[30] : data_i[14];
  assign data_o[15] = head_r ? data_i[31] : data_i[15];
  assign data_o[16] = head_r ? data_i[0] : data_i[16];
  assign data_o[17] = head_r ? data_i[1] : data_i[17];
  assign data_o[18] = head_r ? data_i[2] : data_i[18];
  assign data_o[19] = head_r ? data_i[3] : data_i[19];
  assign data_o[20] = head_r ? data_i[4] : data_i[20];
  assign data_o[21] = head_r ? data_i[5] : data_i[21];
  assign data_o[22] = head_r ? data_i[6] : data_i[22];
  assign data_o[23] = head_r ? data_i[7] : data_i[23];
  assign data_o[24] = head_r ? data_i[8] : data_i[24];
  assign data_o[25] = head_r ? data_i[9] : data_i[25];
  assign data_o[26] = head_r ? data_i[10] : data_i[26];
  assign data_o[27] = head_r ? data_i[11] : data_i[27];
  assign data_o[28] = head_r ? data_i[12] : data_i[28];
  assign data_o[29] = head_r ? data_i[13] : data_i[29];
  assign data_o[30] = head_r ? data_i[14] : data_i[30];
  assign data_o[31] = head_r ? data_i[15] : data_i[31];
  assign v_o[0] = head_r ? v_i[1] : v_i[0];
  assign v_o[1] = head_r ? v_i[0] : v_i[1];
  assign data_o[0] = head_r ? data_i[16] : data_i[0];
  assign data_o[1] = head_r ? data_i[17] : data_i[1];
  assign data_o[2] = head_r ? data_i[18] : data_i[2];
  assign data_o[3] = head_r ? data_i[19] : data_i[3];
  assign data_o[4] = head_r ? data_i[20] : data_i[4];
  assign data_o[5] = head_r ? data_i[21] : data_i[5];
  assign data_o[6] = head_r ? data_i[22] : data_i[6];
  assign data_o[7] = head_r ? data_i[23] : data_i[7];
  assign data_o[8] = head_r ? data_i[24] : data_i[8];
  assign data_o[9] = head_r ? data_i[25] : data_i[9];
  assign data_o[10] = head_r ? data_i[26] : data_i[10];
  always @(posedge clk_i)
    if (reset_i) head_r <= 1'h0;
    else head_r <= _03_;
endmodule
