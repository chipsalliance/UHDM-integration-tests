module bsg_mux(data_i, sel_i, data_o);
  input [15:0] data_i;
  wire [15:0] data_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire \genblk1.unused ;
  input sel_i;
  wire sel_i;
  assign data_o = data_i;
  assign \genblk1.unused  = sel_i;
endmodule
