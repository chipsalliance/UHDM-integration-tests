// We are actually testing including dupliacated packages in Makefile,
// not this module
module top;
endmodule
