module bsg_mux_butterfly(data_i, sel_i, data_o);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  input [511:0] data_i;
  wire [511:0] data_i;
  output [511:0] data_o;
  wire [511:0] data_o;
  wire [3071:0] data_stage;
  wire [31:0] \mux_stage[0].mux_swap[0].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[0].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[0].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[10].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[10].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[10].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[11].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[11].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[11].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[12].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[12].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[12].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[13].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[13].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[13].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[14].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[14].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[14].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[15].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[15].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[15].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[1].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[1].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[1].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[2].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[2].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[2].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[3].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[3].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[3].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[4].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[4].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[4].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[5].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[5].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[5].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[6].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[6].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[6].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[7].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[7].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[7].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[8].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[8].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[8].swap_inst.swap_i ;
  wire [31:0] \mux_stage[0].mux_swap[9].swap_inst.data_i ;
  wire [31:0] \mux_stage[0].mux_swap[9].swap_inst.data_o ;
  wire \mux_stage[0].mux_swap[9].swap_inst.swap_i ;
  wire [63:0] \mux_stage[1].mux_swap[0].swap_inst.data_i ;
  wire [63:0] \mux_stage[1].mux_swap[0].swap_inst.data_o ;
  wire \mux_stage[1].mux_swap[0].swap_inst.swap_i ;
  wire [63:0] \mux_stage[1].mux_swap[1].swap_inst.data_i ;
  wire [63:0] \mux_stage[1].mux_swap[1].swap_inst.data_o ;
  wire \mux_stage[1].mux_swap[1].swap_inst.swap_i ;
  wire [63:0] \mux_stage[1].mux_swap[2].swap_inst.data_i ;
  wire [63:0] \mux_stage[1].mux_swap[2].swap_inst.data_o ;
  wire \mux_stage[1].mux_swap[2].swap_inst.swap_i ;
  wire [63:0] \mux_stage[1].mux_swap[3].swap_inst.data_i ;
  wire [63:0] \mux_stage[1].mux_swap[3].swap_inst.data_o ;
  wire \mux_stage[1].mux_swap[3].swap_inst.swap_i ;
  wire [63:0] \mux_stage[1].mux_swap[4].swap_inst.data_i ;
  wire [63:0] \mux_stage[1].mux_swap[4].swap_inst.data_o ;
  wire \mux_stage[1].mux_swap[4].swap_inst.swap_i ;
  wire [63:0] \mux_stage[1].mux_swap[5].swap_inst.data_i ;
  wire [63:0] \mux_stage[1].mux_swap[5].swap_inst.data_o ;
  wire \mux_stage[1].mux_swap[5].swap_inst.swap_i ;
  wire [63:0] \mux_stage[1].mux_swap[6].swap_inst.data_i ;
  wire [63:0] \mux_stage[1].mux_swap[6].swap_inst.data_o ;
  wire \mux_stage[1].mux_swap[6].swap_inst.swap_i ;
  wire [63:0] \mux_stage[1].mux_swap[7].swap_inst.data_i ;
  wire [63:0] \mux_stage[1].mux_swap[7].swap_inst.data_o ;
  wire \mux_stage[1].mux_swap[7].swap_inst.swap_i ;
  wire [127:0] \mux_stage[2].mux_swap[0].swap_inst.data_i ;
  wire [127:0] \mux_stage[2].mux_swap[0].swap_inst.data_o ;
  wire \mux_stage[2].mux_swap[0].swap_inst.swap_i ;
  wire [127:0] \mux_stage[2].mux_swap[1].swap_inst.data_i ;
  wire [127:0] \mux_stage[2].mux_swap[1].swap_inst.data_o ;
  wire \mux_stage[2].mux_swap[1].swap_inst.swap_i ;
  wire [127:0] \mux_stage[2].mux_swap[2].swap_inst.data_i ;
  wire [127:0] \mux_stage[2].mux_swap[2].swap_inst.data_o ;
  wire \mux_stage[2].mux_swap[2].swap_inst.swap_i ;
  wire [127:0] \mux_stage[2].mux_swap[3].swap_inst.data_i ;
  wire [127:0] \mux_stage[2].mux_swap[3].swap_inst.data_o ;
  wire \mux_stage[2].mux_swap[3].swap_inst.swap_i ;
  wire [255:0] \mux_stage[3].mux_swap[0].swap_inst.data_i ;
  wire [255:0] \mux_stage[3].mux_swap[0].swap_inst.data_o ;
  wire \mux_stage[3].mux_swap[0].swap_inst.swap_i ;
  wire [255:0] \mux_stage[3].mux_swap[1].swap_inst.data_i ;
  wire [255:0] \mux_stage[3].mux_swap[1].swap_inst.data_o ;
  wire \mux_stage[3].mux_swap[1].swap_inst.swap_i ;
  wire [511:0] \mux_stage[4].mux_swap[0].swap_inst.data_i ;
  wire [511:0] \mux_stage[4].mux_swap[0].swap_inst.data_o ;
  wire \mux_stage[4].mux_swap[0].swap_inst.swap_i ;
  input [4:0] sel_i;
  wire [4:0] sel_i;
  assign _0000_ = sel_i[0] ? data_i[16] : data_i[0];
  assign _0001_ = sel_i[0] ? data_i[48] : data_i[32];
  assign _0002_ = sel_i[1] ? _0001_ : _0000_;
  assign _0003_ = sel_i[0] ? data_i[80] : data_i[64];
  assign _0004_ = sel_i[0] ? data_i[112] : data_i[96];
  assign _0005_ = sel_i[1] ? _0004_ : _0003_;
  assign _0006_ = sel_i[2] ? _0005_ : _0002_;
  assign _0007_ = sel_i[0] ? data_i[144] : data_i[128];
  assign _0008_ = sel_i[0] ? data_i[176] : data_i[160];
  assign _0009_ = sel_i[1] ? _0008_ : _0007_;
  assign _0010_ = sel_i[0] ? data_i[208] : data_i[192];
  assign _0011_ = sel_i[0] ? data_i[240] : data_i[224];
  assign _0012_ = sel_i[1] ? _0011_ : _0010_;
  assign _0013_ = sel_i[2] ? _0012_ : _0009_;
  assign _0014_ = sel_i[3] ? _0013_ : _0006_;
  assign _0015_ = sel_i[0] ? data_i[272] : data_i[256];
  assign _0016_ = sel_i[0] ? data_i[304] : data_i[288];
  assign _0017_ = sel_i[1] ? _0016_ : _0015_;
  assign _0018_ = sel_i[0] ? data_i[336] : data_i[320];
  assign _0019_ = sel_i[0] ? data_i[368] : data_i[352];
  assign _0020_ = sel_i[1] ? _0019_ : _0018_;
  assign _0021_ = sel_i[2] ? _0020_ : _0017_;
  assign _0022_ = sel_i[0] ? data_i[400] : data_i[384];
  assign _0023_ = sel_i[0] ? data_i[432] : data_i[416];
  assign _0024_ = sel_i[1] ? _0023_ : _0022_;
  assign _0025_ = sel_i[0] ? data_i[464] : data_i[448];
  assign _0026_ = sel_i[0] ? data_i[496] : data_i[480];
  assign _0027_ = sel_i[1] ? _0026_ : _0025_;
  assign _0028_ = sel_i[2] ? _0027_ : _0024_;
  assign _0029_ = sel_i[3] ? _0028_ : _0021_;
  assign data_o[0] = sel_i[4] ? _0029_ : _0014_;
  assign _0030_ = sel_i[0] ? data_i[17] : data_i[1];
  assign _0031_ = sel_i[0] ? data_i[49] : data_i[33];
  assign _0032_ = sel_i[1] ? _0031_ : _0030_;
  assign _0033_ = sel_i[0] ? data_i[81] : data_i[65];
  assign _0034_ = sel_i[0] ? data_i[113] : data_i[97];
  assign _0035_ = sel_i[1] ? _0034_ : _0033_;
  assign _0036_ = sel_i[2] ? _0035_ : _0032_;
  assign _0037_ = sel_i[0] ? data_i[145] : data_i[129];
  assign _0038_ = sel_i[0] ? data_i[177] : data_i[161];
  assign _0039_ = sel_i[1] ? _0038_ : _0037_;
  assign _0040_ = sel_i[0] ? data_i[209] : data_i[193];
  assign _0041_ = sel_i[0] ? data_i[241] : data_i[225];
  assign _0042_ = sel_i[1] ? _0041_ : _0040_;
  assign _0043_ = sel_i[2] ? _0042_ : _0039_;
  assign _0044_ = sel_i[3] ? _0043_ : _0036_;
  assign _0045_ = sel_i[0] ? data_i[273] : data_i[257];
  assign _0046_ = sel_i[0] ? data_i[305] : data_i[289];
  assign _0047_ = sel_i[1] ? _0046_ : _0045_;
  assign _0048_ = sel_i[0] ? data_i[337] : data_i[321];
  assign _0049_ = sel_i[0] ? data_i[369] : data_i[353];
  assign _0050_ = sel_i[1] ? _0049_ : _0048_;
  assign _0051_ = sel_i[2] ? _0050_ : _0047_;
  assign _0052_ = sel_i[0] ? data_i[401] : data_i[385];
  assign _0053_ = sel_i[0] ? data_i[433] : data_i[417];
  assign _0054_ = sel_i[1] ? _0053_ : _0052_;
  assign _0055_ = sel_i[0] ? data_i[465] : data_i[449];
  assign _0056_ = sel_i[0] ? data_i[497] : data_i[481];
  assign _0057_ = sel_i[1] ? _0056_ : _0055_;
  assign _0058_ = sel_i[2] ? _0057_ : _0054_;
  assign _0059_ = sel_i[3] ? _0058_ : _0051_;
  assign data_o[1] = sel_i[4] ? _0059_ : _0044_;
  assign _0060_ = sel_i[0] ? data_i[18] : data_i[2];
  assign _0061_ = sel_i[0] ? data_i[50] : data_i[34];
  assign _0062_ = sel_i[1] ? _0061_ : _0060_;
  assign _0063_ = sel_i[0] ? data_i[82] : data_i[66];
  assign _0064_ = sel_i[0] ? data_i[114] : data_i[98];
  assign _0065_ = sel_i[1] ? _0064_ : _0063_;
  assign _0066_ = sel_i[2] ? _0065_ : _0062_;
  assign _0067_ = sel_i[0] ? data_i[146] : data_i[130];
  assign _0068_ = sel_i[0] ? data_i[178] : data_i[162];
  assign _0069_ = sel_i[1] ? _0068_ : _0067_;
  assign _0070_ = sel_i[0] ? data_i[210] : data_i[194];
  assign _0071_ = sel_i[0] ? data_i[242] : data_i[226];
  assign _0072_ = sel_i[1] ? _0071_ : _0070_;
  assign _0073_ = sel_i[2] ? _0072_ : _0069_;
  assign _0074_ = sel_i[3] ? _0073_ : _0066_;
  assign _0075_ = sel_i[0] ? data_i[274] : data_i[258];
  assign _0076_ = sel_i[0] ? data_i[306] : data_i[290];
  assign _0077_ = sel_i[1] ? _0076_ : _0075_;
  assign _0078_ = sel_i[0] ? data_i[338] : data_i[322];
  assign _0079_ = sel_i[0] ? data_i[370] : data_i[354];
  assign _0080_ = sel_i[1] ? _0079_ : _0078_;
  assign _0081_ = sel_i[2] ? _0080_ : _0077_;
  assign _0082_ = sel_i[0] ? data_i[402] : data_i[386];
  assign _0083_ = sel_i[0] ? data_i[434] : data_i[418];
  assign _0084_ = sel_i[1] ? _0083_ : _0082_;
  assign _0085_ = sel_i[0] ? data_i[466] : data_i[450];
  assign _0086_ = sel_i[0] ? data_i[498] : data_i[482];
  assign _0087_ = sel_i[1] ? _0086_ : _0085_;
  assign _0088_ = sel_i[2] ? _0087_ : _0084_;
  assign _0089_ = sel_i[3] ? _0088_ : _0081_;
  assign data_o[2] = sel_i[4] ? _0089_ : _0074_;
  assign _0090_ = sel_i[0] ? data_i[19] : data_i[3];
  assign _0091_ = sel_i[0] ? data_i[51] : data_i[35];
  assign _0092_ = sel_i[1] ? _0091_ : _0090_;
  assign _0093_ = sel_i[0] ? data_i[83] : data_i[67];
  assign _0094_ = sel_i[0] ? data_i[115] : data_i[99];
  assign _0095_ = sel_i[1] ? _0094_ : _0093_;
  assign _0096_ = sel_i[2] ? _0095_ : _0092_;
  assign _0097_ = sel_i[0] ? data_i[147] : data_i[131];
  assign _0098_ = sel_i[0] ? data_i[179] : data_i[163];
  assign _0099_ = sel_i[1] ? _0098_ : _0097_;
  assign _0100_ = sel_i[0] ? data_i[211] : data_i[195];
  assign _0101_ = sel_i[0] ? data_i[243] : data_i[227];
  assign _0102_ = sel_i[1] ? _0101_ : _0100_;
  assign _0103_ = sel_i[2] ? _0102_ : _0099_;
  assign _0104_ = sel_i[3] ? _0103_ : _0096_;
  assign _0105_ = sel_i[0] ? data_i[275] : data_i[259];
  assign _0106_ = sel_i[0] ? data_i[307] : data_i[291];
  assign _0107_ = sel_i[1] ? _0106_ : _0105_;
  assign _0108_ = sel_i[0] ? data_i[339] : data_i[323];
  assign _0109_ = sel_i[0] ? data_i[371] : data_i[355];
  assign _0110_ = sel_i[1] ? _0109_ : _0108_;
  assign _0111_ = sel_i[2] ? _0110_ : _0107_;
  assign _0112_ = sel_i[0] ? data_i[403] : data_i[387];
  assign _0113_ = sel_i[0] ? data_i[435] : data_i[419];
  assign _0114_ = sel_i[1] ? _0113_ : _0112_;
  assign _0115_ = sel_i[0] ? data_i[467] : data_i[451];
  assign _0116_ = sel_i[0] ? data_i[499] : data_i[483];
  assign _0117_ = sel_i[1] ? _0116_ : _0115_;
  assign _0118_ = sel_i[2] ? _0117_ : _0114_;
  assign _0119_ = sel_i[3] ? _0118_ : _0111_;
  assign data_o[3] = sel_i[4] ? _0119_ : _0104_;
  assign _0120_ = sel_i[0] ? data_i[20] : data_i[4];
  assign _0121_ = sel_i[0] ? data_i[52] : data_i[36];
  assign _0122_ = sel_i[1] ? _0121_ : _0120_;
  assign _0123_ = sel_i[0] ? data_i[84] : data_i[68];
  assign _0124_ = sel_i[0] ? data_i[116] : data_i[100];
  assign _0125_ = sel_i[1] ? _0124_ : _0123_;
  assign _0126_ = sel_i[2] ? _0125_ : _0122_;
  assign _0127_ = sel_i[0] ? data_i[148] : data_i[132];
  assign _0128_ = sel_i[0] ? data_i[180] : data_i[164];
  assign _0129_ = sel_i[1] ? _0128_ : _0127_;
  assign _0130_ = sel_i[0] ? data_i[212] : data_i[196];
  assign _0131_ = sel_i[0] ? data_i[244] : data_i[228];
  assign _0132_ = sel_i[1] ? _0131_ : _0130_;
  assign _0133_ = sel_i[2] ? _0132_ : _0129_;
  assign _0134_ = sel_i[3] ? _0133_ : _0126_;
  assign _0135_ = sel_i[0] ? data_i[276] : data_i[260];
  assign _0136_ = sel_i[0] ? data_i[308] : data_i[292];
  assign _0137_ = sel_i[1] ? _0136_ : _0135_;
  assign _0138_ = sel_i[0] ? data_i[340] : data_i[324];
  assign _0139_ = sel_i[0] ? data_i[372] : data_i[356];
  assign _0140_ = sel_i[1] ? _0139_ : _0138_;
  assign _0141_ = sel_i[2] ? _0140_ : _0137_;
  assign _0142_ = sel_i[0] ? data_i[404] : data_i[388];
  assign _0143_ = sel_i[0] ? data_i[436] : data_i[420];
  assign _0144_ = sel_i[1] ? _0143_ : _0142_;
  assign _0145_ = sel_i[0] ? data_i[468] : data_i[452];
  assign _0146_ = sel_i[0] ? data_i[500] : data_i[484];
  assign _0147_ = sel_i[1] ? _0146_ : _0145_;
  assign _0148_ = sel_i[2] ? _0147_ : _0144_;
  assign _0149_ = sel_i[3] ? _0148_ : _0141_;
  assign data_o[4] = sel_i[4] ? _0149_ : _0134_;
  assign _0150_ = sel_i[0] ? data_i[21] : data_i[5];
  assign _0151_ = sel_i[0] ? data_i[53] : data_i[37];
  assign _0152_ = sel_i[1] ? _0151_ : _0150_;
  assign _0153_ = sel_i[0] ? data_i[85] : data_i[69];
  assign _0154_ = sel_i[0] ? data_i[117] : data_i[101];
  assign _0155_ = sel_i[1] ? _0154_ : _0153_;
  assign _0156_ = sel_i[2] ? _0155_ : _0152_;
  assign _0157_ = sel_i[0] ? data_i[149] : data_i[133];
  assign _0158_ = sel_i[0] ? data_i[181] : data_i[165];
  assign _0159_ = sel_i[1] ? _0158_ : _0157_;
  assign _0160_ = sel_i[0] ? data_i[213] : data_i[197];
  assign _0161_ = sel_i[0] ? data_i[245] : data_i[229];
  assign _0162_ = sel_i[1] ? _0161_ : _0160_;
  assign _0163_ = sel_i[2] ? _0162_ : _0159_;
  assign _0164_ = sel_i[3] ? _0163_ : _0156_;
  assign _0165_ = sel_i[0] ? data_i[277] : data_i[261];
  assign _0166_ = sel_i[0] ? data_i[309] : data_i[293];
  assign _0167_ = sel_i[1] ? _0166_ : _0165_;
  assign _0168_ = sel_i[0] ? data_i[341] : data_i[325];
  assign _0169_ = sel_i[0] ? data_i[373] : data_i[357];
  assign _0170_ = sel_i[1] ? _0169_ : _0168_;
  assign _0171_ = sel_i[2] ? _0170_ : _0167_;
  assign _0172_ = sel_i[0] ? data_i[405] : data_i[389];
  assign _0173_ = sel_i[0] ? data_i[437] : data_i[421];
  assign _0174_ = sel_i[1] ? _0173_ : _0172_;
  assign _0175_ = sel_i[0] ? data_i[469] : data_i[453];
  assign _0176_ = sel_i[0] ? data_i[501] : data_i[485];
  assign _0177_ = sel_i[1] ? _0176_ : _0175_;
  assign _0178_ = sel_i[2] ? _0177_ : _0174_;
  assign _0179_ = sel_i[3] ? _0178_ : _0171_;
  assign data_o[5] = sel_i[4] ? _0179_ : _0164_;
  assign _0180_ = sel_i[0] ? data_i[22] : data_i[6];
  assign _0181_ = sel_i[0] ? data_i[54] : data_i[38];
  assign _0182_ = sel_i[1] ? _0181_ : _0180_;
  assign _0183_ = sel_i[0] ? data_i[86] : data_i[70];
  assign _0184_ = sel_i[0] ? data_i[118] : data_i[102];
  assign _0185_ = sel_i[1] ? _0184_ : _0183_;
  assign _0186_ = sel_i[2] ? _0185_ : _0182_;
  assign _0187_ = sel_i[0] ? data_i[150] : data_i[134];
  assign _0188_ = sel_i[0] ? data_i[182] : data_i[166];
  assign _0189_ = sel_i[1] ? _0188_ : _0187_;
  assign _0190_ = sel_i[0] ? data_i[214] : data_i[198];
  assign _0191_ = sel_i[0] ? data_i[246] : data_i[230];
  assign _0192_ = sel_i[1] ? _0191_ : _0190_;
  assign _0193_ = sel_i[2] ? _0192_ : _0189_;
  assign _0194_ = sel_i[3] ? _0193_ : _0186_;
  assign _0195_ = sel_i[0] ? data_i[278] : data_i[262];
  assign _0196_ = sel_i[0] ? data_i[310] : data_i[294];
  assign _0197_ = sel_i[1] ? _0196_ : _0195_;
  assign _0198_ = sel_i[0] ? data_i[342] : data_i[326];
  assign _0199_ = sel_i[0] ? data_i[374] : data_i[358];
  assign _0200_ = sel_i[1] ? _0199_ : _0198_;
  assign _0201_ = sel_i[2] ? _0200_ : _0197_;
  assign _0202_ = sel_i[0] ? data_i[406] : data_i[390];
  assign _0203_ = sel_i[0] ? data_i[438] : data_i[422];
  assign _0204_ = sel_i[1] ? _0203_ : _0202_;
  assign _0205_ = sel_i[0] ? data_i[470] : data_i[454];
  assign _0206_ = sel_i[0] ? data_i[502] : data_i[486];
  assign _0207_ = sel_i[1] ? _0206_ : _0205_;
  assign _0208_ = sel_i[2] ? _0207_ : _0204_;
  assign _0209_ = sel_i[3] ? _0208_ : _0201_;
  assign data_o[6] = sel_i[4] ? _0209_ : _0194_;
  assign _0210_ = sel_i[0] ? data_i[23] : data_i[7];
  assign _0211_ = sel_i[0] ? data_i[55] : data_i[39];
  assign _0212_ = sel_i[1] ? _0211_ : _0210_;
  assign _0213_ = sel_i[0] ? data_i[87] : data_i[71];
  assign _0214_ = sel_i[0] ? data_i[119] : data_i[103];
  assign _0215_ = sel_i[1] ? _0214_ : _0213_;
  assign _0216_ = sel_i[2] ? _0215_ : _0212_;
  assign _0217_ = sel_i[0] ? data_i[151] : data_i[135];
  assign _0218_ = sel_i[0] ? data_i[183] : data_i[167];
  assign _0219_ = sel_i[1] ? _0218_ : _0217_;
  assign _0220_ = sel_i[0] ? data_i[215] : data_i[199];
  assign _0221_ = sel_i[0] ? data_i[247] : data_i[231];
  assign _0222_ = sel_i[1] ? _0221_ : _0220_;
  assign _0223_ = sel_i[2] ? _0222_ : _0219_;
  assign _0224_ = sel_i[3] ? _0223_ : _0216_;
  assign _0225_ = sel_i[0] ? data_i[279] : data_i[263];
  assign _0226_ = sel_i[0] ? data_i[311] : data_i[295];
  assign _0227_ = sel_i[1] ? _0226_ : _0225_;
  assign _0228_ = sel_i[0] ? data_i[343] : data_i[327];
  assign _0229_ = sel_i[0] ? data_i[375] : data_i[359];
  assign _0230_ = sel_i[1] ? _0229_ : _0228_;
  assign _0231_ = sel_i[2] ? _0230_ : _0227_;
  assign _0232_ = sel_i[0] ? data_i[407] : data_i[391];
  assign _0233_ = sel_i[0] ? data_i[439] : data_i[423];
  assign _0234_ = sel_i[1] ? _0233_ : _0232_;
  assign _0235_ = sel_i[0] ? data_i[471] : data_i[455];
  assign _0236_ = sel_i[0] ? data_i[503] : data_i[487];
  assign _0237_ = sel_i[1] ? _0236_ : _0235_;
  assign _0238_ = sel_i[2] ? _0237_ : _0234_;
  assign _0239_ = sel_i[3] ? _0238_ : _0231_;
  assign data_o[7] = sel_i[4] ? _0239_ : _0224_;
  assign _0240_ = sel_i[0] ? data_i[24] : data_i[8];
  assign _0241_ = sel_i[0] ? data_i[56] : data_i[40];
  assign _0242_ = sel_i[1] ? _0241_ : _0240_;
  assign _0243_ = sel_i[0] ? data_i[88] : data_i[72];
  assign _0244_ = sel_i[0] ? data_i[120] : data_i[104];
  assign _0245_ = sel_i[1] ? _0244_ : _0243_;
  assign _0246_ = sel_i[2] ? _0245_ : _0242_;
  assign _0247_ = sel_i[0] ? data_i[152] : data_i[136];
  assign _0248_ = sel_i[0] ? data_i[184] : data_i[168];
  assign _0249_ = sel_i[1] ? _0248_ : _0247_;
  assign _0250_ = sel_i[0] ? data_i[216] : data_i[200];
  assign _0251_ = sel_i[0] ? data_i[248] : data_i[232];
  assign _0252_ = sel_i[1] ? _0251_ : _0250_;
  assign _0253_ = sel_i[2] ? _0252_ : _0249_;
  assign _0254_ = sel_i[3] ? _0253_ : _0246_;
  assign _0255_ = sel_i[0] ? data_i[280] : data_i[264];
  assign _0256_ = sel_i[0] ? data_i[312] : data_i[296];
  assign _0257_ = sel_i[1] ? _0256_ : _0255_;
  assign _0258_ = sel_i[0] ? data_i[344] : data_i[328];
  assign _0259_ = sel_i[0] ? data_i[376] : data_i[360];
  assign _0260_ = sel_i[1] ? _0259_ : _0258_;
  assign _0261_ = sel_i[2] ? _0260_ : _0257_;
  assign _0262_ = sel_i[0] ? data_i[408] : data_i[392];
  assign _0263_ = sel_i[0] ? data_i[440] : data_i[424];
  assign _0264_ = sel_i[1] ? _0263_ : _0262_;
  assign _0265_ = sel_i[0] ? data_i[472] : data_i[456];
  assign _0266_ = sel_i[0] ? data_i[504] : data_i[488];
  assign _0267_ = sel_i[1] ? _0266_ : _0265_;
  assign _0268_ = sel_i[2] ? _0267_ : _0264_;
  assign _0269_ = sel_i[3] ? _0268_ : _0261_;
  assign data_o[8] = sel_i[4] ? _0269_ : _0254_;
  assign _0270_ = sel_i[0] ? data_i[25] : data_i[9];
  assign _0271_ = sel_i[0] ? data_i[57] : data_i[41];
  assign _0272_ = sel_i[1] ? _0271_ : _0270_;
  assign _0273_ = sel_i[0] ? data_i[89] : data_i[73];
  assign _0274_ = sel_i[0] ? data_i[121] : data_i[105];
  assign _0275_ = sel_i[1] ? _0274_ : _0273_;
  assign _0276_ = sel_i[2] ? _0275_ : _0272_;
  assign _0277_ = sel_i[0] ? data_i[153] : data_i[137];
  assign _0278_ = sel_i[0] ? data_i[185] : data_i[169];
  assign _0279_ = sel_i[1] ? _0278_ : _0277_;
  assign _0280_ = sel_i[0] ? data_i[217] : data_i[201];
  assign _0281_ = sel_i[0] ? data_i[249] : data_i[233];
  assign _0282_ = sel_i[1] ? _0281_ : _0280_;
  assign _0283_ = sel_i[2] ? _0282_ : _0279_;
  assign _0284_ = sel_i[3] ? _0283_ : _0276_;
  assign _0285_ = sel_i[0] ? data_i[281] : data_i[265];
  assign _0286_ = sel_i[0] ? data_i[313] : data_i[297];
  assign _0287_ = sel_i[1] ? _0286_ : _0285_;
  assign _0288_ = sel_i[0] ? data_i[345] : data_i[329];
  assign _0289_ = sel_i[0] ? data_i[377] : data_i[361];
  assign _0290_ = sel_i[1] ? _0289_ : _0288_;
  assign _0291_ = sel_i[2] ? _0290_ : _0287_;
  assign _0292_ = sel_i[0] ? data_i[409] : data_i[393];
  assign _0293_ = sel_i[0] ? data_i[441] : data_i[425];
  assign _0294_ = sel_i[1] ? _0293_ : _0292_;
  assign _0295_ = sel_i[0] ? data_i[473] : data_i[457];
  assign _0296_ = sel_i[0] ? data_i[505] : data_i[489];
  assign _0297_ = sel_i[1] ? _0296_ : _0295_;
  assign _0298_ = sel_i[2] ? _0297_ : _0294_;
  assign _0299_ = sel_i[3] ? _0298_ : _0291_;
  assign data_o[9] = sel_i[4] ? _0299_ : _0284_;
  assign _0300_ = sel_i[0] ? data_i[26] : data_i[10];
  assign _0301_ = sel_i[0] ? data_i[58] : data_i[42];
  assign _0302_ = sel_i[1] ? _0301_ : _0300_;
  assign _0303_ = sel_i[0] ? data_i[90] : data_i[74];
  assign _0304_ = sel_i[0] ? data_i[122] : data_i[106];
  assign _0305_ = sel_i[1] ? _0304_ : _0303_;
  assign _0306_ = sel_i[2] ? _0305_ : _0302_;
  assign _0307_ = sel_i[0] ? data_i[154] : data_i[138];
  assign _0308_ = sel_i[0] ? data_i[186] : data_i[170];
  assign _0309_ = sel_i[1] ? _0308_ : _0307_;
  assign _0310_ = sel_i[0] ? data_i[218] : data_i[202];
  assign _0311_ = sel_i[0] ? data_i[250] : data_i[234];
  assign _0312_ = sel_i[1] ? _0311_ : _0310_;
  assign _0313_ = sel_i[2] ? _0312_ : _0309_;
  assign _0314_ = sel_i[3] ? _0313_ : _0306_;
  assign _0315_ = sel_i[0] ? data_i[282] : data_i[266];
  assign _0316_ = sel_i[0] ? data_i[314] : data_i[298];
  assign _0317_ = sel_i[1] ? _0316_ : _0315_;
  assign _0318_ = sel_i[0] ? data_i[346] : data_i[330];
  assign _0319_ = sel_i[0] ? data_i[378] : data_i[362];
  assign _0320_ = sel_i[1] ? _0319_ : _0318_;
  assign _0321_ = sel_i[2] ? _0320_ : _0317_;
  assign _0322_ = sel_i[0] ? data_i[410] : data_i[394];
  assign _0323_ = sel_i[0] ? data_i[442] : data_i[426];
  assign _0324_ = sel_i[1] ? _0323_ : _0322_;
  assign _0325_ = sel_i[0] ? data_i[474] : data_i[458];
  assign _0326_ = sel_i[0] ? data_i[506] : data_i[490];
  assign _0327_ = sel_i[1] ? _0326_ : _0325_;
  assign _0328_ = sel_i[2] ? _0327_ : _0324_;
  assign _0329_ = sel_i[3] ? _0328_ : _0321_;
  assign data_o[10] = sel_i[4] ? _0329_ : _0314_;
  assign _0330_ = sel_i[0] ? data_i[27] : data_i[11];
  assign _0331_ = sel_i[0] ? data_i[59] : data_i[43];
  assign _0332_ = sel_i[1] ? _0331_ : _0330_;
  assign _0333_ = sel_i[0] ? data_i[91] : data_i[75];
  assign _0334_ = sel_i[0] ? data_i[123] : data_i[107];
  assign _0335_ = sel_i[1] ? _0334_ : _0333_;
  assign _0336_ = sel_i[2] ? _0335_ : _0332_;
  assign _0337_ = sel_i[0] ? data_i[155] : data_i[139];
  assign _0338_ = sel_i[0] ? data_i[187] : data_i[171];
  assign _0339_ = sel_i[1] ? _0338_ : _0337_;
  assign _0340_ = sel_i[0] ? data_i[219] : data_i[203];
  assign _0341_ = sel_i[0] ? data_i[251] : data_i[235];
  assign _0342_ = sel_i[1] ? _0341_ : _0340_;
  assign _0343_ = sel_i[2] ? _0342_ : _0339_;
  assign _0344_ = sel_i[3] ? _0343_ : _0336_;
  assign _0345_ = sel_i[0] ? data_i[283] : data_i[267];
  assign _0346_ = sel_i[0] ? data_i[315] : data_i[299];
  assign _0347_ = sel_i[1] ? _0346_ : _0345_;
  assign _0348_ = sel_i[0] ? data_i[347] : data_i[331];
  assign _0349_ = sel_i[0] ? data_i[379] : data_i[363];
  assign _0350_ = sel_i[1] ? _0349_ : _0348_;
  assign _0351_ = sel_i[2] ? _0350_ : _0347_;
  assign _0352_ = sel_i[0] ? data_i[411] : data_i[395];
  assign _0353_ = sel_i[0] ? data_i[443] : data_i[427];
  assign _0354_ = sel_i[1] ? _0353_ : _0352_;
  assign _0355_ = sel_i[0] ? data_i[475] : data_i[459];
  assign _0356_ = sel_i[0] ? data_i[507] : data_i[491];
  assign _0357_ = sel_i[1] ? _0356_ : _0355_;
  assign _0358_ = sel_i[2] ? _0357_ : _0354_;
  assign _0359_ = sel_i[3] ? _0358_ : _0351_;
  assign data_o[11] = sel_i[4] ? _0359_ : _0344_;
  assign _0360_ = sel_i[0] ? data_i[28] : data_i[12];
  assign _0361_ = sel_i[0] ? data_i[60] : data_i[44];
  assign _0362_ = sel_i[1] ? _0361_ : _0360_;
  assign _0363_ = sel_i[0] ? data_i[92] : data_i[76];
  assign _0364_ = sel_i[0] ? data_i[124] : data_i[108];
  assign _0365_ = sel_i[1] ? _0364_ : _0363_;
  assign _0366_ = sel_i[2] ? _0365_ : _0362_;
  assign _0367_ = sel_i[0] ? data_i[156] : data_i[140];
  assign _0368_ = sel_i[0] ? data_i[188] : data_i[172];
  assign _0369_ = sel_i[1] ? _0368_ : _0367_;
  assign _0370_ = sel_i[0] ? data_i[220] : data_i[204];
  assign _0371_ = sel_i[0] ? data_i[252] : data_i[236];
  assign _0372_ = sel_i[1] ? _0371_ : _0370_;
  assign _0373_ = sel_i[2] ? _0372_ : _0369_;
  assign _0374_ = sel_i[3] ? _0373_ : _0366_;
  assign _0375_ = sel_i[0] ? data_i[284] : data_i[268];
  assign _0376_ = sel_i[0] ? data_i[316] : data_i[300];
  assign _0377_ = sel_i[1] ? _0376_ : _0375_;
  assign _0378_ = sel_i[0] ? data_i[348] : data_i[332];
  assign _0379_ = sel_i[0] ? data_i[380] : data_i[364];
  assign _0380_ = sel_i[1] ? _0379_ : _0378_;
  assign _0381_ = sel_i[2] ? _0380_ : _0377_;
  assign _0382_ = sel_i[0] ? data_i[412] : data_i[396];
  assign _0383_ = sel_i[0] ? data_i[444] : data_i[428];
  assign _0384_ = sel_i[1] ? _0383_ : _0382_;
  assign _0385_ = sel_i[0] ? data_i[476] : data_i[460];
  assign _0386_ = sel_i[0] ? data_i[508] : data_i[492];
  assign _0387_ = sel_i[1] ? _0386_ : _0385_;
  assign _0388_ = sel_i[2] ? _0387_ : _0384_;
  assign _0389_ = sel_i[3] ? _0388_ : _0381_;
  assign data_o[12] = sel_i[4] ? _0389_ : _0374_;
  assign _0390_ = sel_i[0] ? data_i[29] : data_i[13];
  assign _0391_ = sel_i[0] ? data_i[61] : data_i[45];
  assign _0392_ = sel_i[1] ? _0391_ : _0390_;
  assign _0393_ = sel_i[0] ? data_i[93] : data_i[77];
  assign _0394_ = sel_i[0] ? data_i[125] : data_i[109];
  assign _0395_ = sel_i[1] ? _0394_ : _0393_;
  assign _0396_ = sel_i[2] ? _0395_ : _0392_;
  assign _0397_ = sel_i[0] ? data_i[157] : data_i[141];
  assign _0398_ = sel_i[0] ? data_i[189] : data_i[173];
  assign _0399_ = sel_i[1] ? _0398_ : _0397_;
  assign _0400_ = sel_i[0] ? data_i[221] : data_i[205];
  assign _0401_ = sel_i[0] ? data_i[253] : data_i[237];
  assign _0402_ = sel_i[1] ? _0401_ : _0400_;
  assign _0403_ = sel_i[2] ? _0402_ : _0399_;
  assign _0404_ = sel_i[3] ? _0403_ : _0396_;
  assign _0405_ = sel_i[0] ? data_i[285] : data_i[269];
  assign _0406_ = sel_i[0] ? data_i[317] : data_i[301];
  assign _0407_ = sel_i[1] ? _0406_ : _0405_;
  assign _0408_ = sel_i[0] ? data_i[349] : data_i[333];
  assign _0409_ = sel_i[0] ? data_i[381] : data_i[365];
  assign _0410_ = sel_i[1] ? _0409_ : _0408_;
  assign _0411_ = sel_i[2] ? _0410_ : _0407_;
  assign _0412_ = sel_i[0] ? data_i[413] : data_i[397];
  assign _0413_ = sel_i[0] ? data_i[445] : data_i[429];
  assign _0414_ = sel_i[1] ? _0413_ : _0412_;
  assign _0415_ = sel_i[0] ? data_i[477] : data_i[461];
  assign _0416_ = sel_i[0] ? data_i[509] : data_i[493];
  assign _0417_ = sel_i[1] ? _0416_ : _0415_;
  assign _0418_ = sel_i[2] ? _0417_ : _0414_;
  assign _0419_ = sel_i[3] ? _0418_ : _0411_;
  assign data_o[13] = sel_i[4] ? _0419_ : _0404_;
  assign _0420_ = sel_i[0] ? data_i[30] : data_i[14];
  assign _0421_ = sel_i[0] ? data_i[62] : data_i[46];
  assign _0422_ = sel_i[1] ? _0421_ : _0420_;
  assign _0423_ = sel_i[0] ? data_i[94] : data_i[78];
  assign _0424_ = sel_i[0] ? data_i[126] : data_i[110];
  assign _0425_ = sel_i[1] ? _0424_ : _0423_;
  assign _0426_ = sel_i[2] ? _0425_ : _0422_;
  assign _0427_ = sel_i[0] ? data_i[158] : data_i[142];
  assign _0428_ = sel_i[0] ? data_i[190] : data_i[174];
  assign _0429_ = sel_i[1] ? _0428_ : _0427_;
  assign _0430_ = sel_i[0] ? data_i[222] : data_i[206];
  assign _0431_ = sel_i[0] ? data_i[254] : data_i[238];
  assign _0432_ = sel_i[1] ? _0431_ : _0430_;
  assign _0433_ = sel_i[2] ? _0432_ : _0429_;
  assign _0434_ = sel_i[3] ? _0433_ : _0426_;
  assign _0435_ = sel_i[0] ? data_i[286] : data_i[270];
  assign _0436_ = sel_i[0] ? data_i[318] : data_i[302];
  assign _0437_ = sel_i[1] ? _0436_ : _0435_;
  assign _0438_ = sel_i[0] ? data_i[350] : data_i[334];
  assign _0439_ = sel_i[0] ? data_i[382] : data_i[366];
  assign _0440_ = sel_i[1] ? _0439_ : _0438_;
  assign _0441_ = sel_i[2] ? _0440_ : _0437_;
  assign _0442_ = sel_i[0] ? data_i[414] : data_i[398];
  assign _0443_ = sel_i[0] ? data_i[446] : data_i[430];
  assign _0444_ = sel_i[1] ? _0443_ : _0442_;
  assign _0445_ = sel_i[0] ? data_i[478] : data_i[462];
  assign _0446_ = sel_i[0] ? data_i[510] : data_i[494];
  assign _0447_ = sel_i[1] ? _0446_ : _0445_;
  assign _0448_ = sel_i[2] ? _0447_ : _0444_;
  assign _0449_ = sel_i[3] ? _0448_ : _0441_;
  assign data_o[14] = sel_i[4] ? _0449_ : _0434_;
  assign _0450_ = sel_i[0] ? data_i[31] : data_i[15];
  assign _0451_ = sel_i[0] ? data_i[63] : data_i[47];
  assign _0452_ = sel_i[1] ? _0451_ : _0450_;
  assign _0453_ = sel_i[0] ? data_i[95] : data_i[79];
  assign _0454_ = sel_i[0] ? data_i[127] : data_i[111];
  assign _0455_ = sel_i[1] ? _0454_ : _0453_;
  assign _0456_ = sel_i[2] ? _0455_ : _0452_;
  assign _0457_ = sel_i[0] ? data_i[159] : data_i[143];
  assign _0458_ = sel_i[0] ? data_i[191] : data_i[175];
  assign _0459_ = sel_i[1] ? _0458_ : _0457_;
  assign _0460_ = sel_i[0] ? data_i[223] : data_i[207];
  assign _0461_ = sel_i[0] ? data_i[255] : data_i[239];
  assign _0462_ = sel_i[1] ? _0461_ : _0460_;
  assign _0463_ = sel_i[2] ? _0462_ : _0459_;
  assign _0464_ = sel_i[3] ? _0463_ : _0456_;
  assign _0465_ = sel_i[0] ? data_i[287] : data_i[271];
  assign _0466_ = sel_i[0] ? data_i[319] : data_i[303];
  assign _0467_ = sel_i[1] ? _0466_ : _0465_;
  assign _0468_ = sel_i[0] ? data_i[351] : data_i[335];
  assign _0469_ = sel_i[0] ? data_i[383] : data_i[367];
  assign _0470_ = sel_i[1] ? _0469_ : _0468_;
  assign _0471_ = sel_i[2] ? _0470_ : _0467_;
  assign _0472_ = sel_i[0] ? data_i[415] : data_i[399];
  assign _0473_ = sel_i[0] ? data_i[447] : data_i[431];
  assign _0474_ = sel_i[1] ? _0473_ : _0472_;
  assign _0475_ = sel_i[0] ? data_i[479] : data_i[463];
  assign _0476_ = sel_i[0] ? data_i[511] : data_i[495];
  assign _0477_ = sel_i[1] ? _0476_ : _0475_;
  assign _0478_ = sel_i[2] ? _0477_ : _0474_;
  assign _0479_ = sel_i[3] ? _0478_ : _0471_;
  assign data_o[15] = sel_i[4] ? _0479_ : _0464_;
  assign _0480_ = sel_i[0] ? data_i[0] : data_i[16];
  assign _0481_ = sel_i[0] ? data_i[32] : data_i[48];
  assign _0482_ = sel_i[1] ? _0481_ : _0480_;
  assign _0483_ = sel_i[0] ? data_i[64] : data_i[80];
  assign _0484_ = sel_i[0] ? data_i[96] : data_i[112];
  assign _0485_ = sel_i[1] ? _0484_ : _0483_;
  assign _0486_ = sel_i[2] ? _0485_ : _0482_;
  assign _0487_ = sel_i[0] ? data_i[128] : data_i[144];
  assign _0488_ = sel_i[0] ? data_i[160] : data_i[176];
  assign _0489_ = sel_i[1] ? _0488_ : _0487_;
  assign _0490_ = sel_i[0] ? data_i[192] : data_i[208];
  assign _0491_ = sel_i[0] ? data_i[224] : data_i[240];
  assign _0492_ = sel_i[1] ? _0491_ : _0490_;
  assign _0493_ = sel_i[2] ? _0492_ : _0489_;
  assign _0494_ = sel_i[3] ? _0493_ : _0486_;
  assign _0495_ = sel_i[0] ? data_i[256] : data_i[272];
  assign _0496_ = sel_i[0] ? data_i[288] : data_i[304];
  assign _0497_ = sel_i[1] ? _0496_ : _0495_;
  assign _0498_ = sel_i[0] ? data_i[320] : data_i[336];
  assign _0499_ = sel_i[0] ? data_i[352] : data_i[368];
  assign _0500_ = sel_i[1] ? _0499_ : _0498_;
  assign _0501_ = sel_i[2] ? _0500_ : _0497_;
  assign _0502_ = sel_i[0] ? data_i[384] : data_i[400];
  assign _0503_ = sel_i[0] ? data_i[416] : data_i[432];
  assign _0504_ = sel_i[1] ? _0503_ : _0502_;
  assign _0505_ = sel_i[0] ? data_i[448] : data_i[464];
  assign _0506_ = sel_i[0] ? data_i[480] : data_i[496];
  assign _0507_ = sel_i[1] ? _0506_ : _0505_;
  assign _0508_ = sel_i[2] ? _0507_ : _0504_;
  assign _0509_ = sel_i[3] ? _0508_ : _0501_;
  assign data_o[16] = sel_i[4] ? _0509_ : _0494_;
  assign _0510_ = sel_i[0] ? data_i[1] : data_i[17];
  assign _0511_ = sel_i[0] ? data_i[33] : data_i[49];
  assign _0512_ = sel_i[1] ? _0511_ : _0510_;
  assign _0513_ = sel_i[0] ? data_i[65] : data_i[81];
  assign _0514_ = sel_i[0] ? data_i[97] : data_i[113];
  assign _0515_ = sel_i[1] ? _0514_ : _0513_;
  assign _0516_ = sel_i[2] ? _0515_ : _0512_;
  assign _0517_ = sel_i[0] ? data_i[129] : data_i[145];
  assign _0518_ = sel_i[0] ? data_i[161] : data_i[177];
  assign _0519_ = sel_i[1] ? _0518_ : _0517_;
  assign _0520_ = sel_i[0] ? data_i[193] : data_i[209];
  assign _0521_ = sel_i[0] ? data_i[225] : data_i[241];
  assign _0522_ = sel_i[1] ? _0521_ : _0520_;
  assign _0523_ = sel_i[2] ? _0522_ : _0519_;
  assign _0524_ = sel_i[3] ? _0523_ : _0516_;
  assign _0525_ = sel_i[0] ? data_i[257] : data_i[273];
  assign _0526_ = sel_i[0] ? data_i[289] : data_i[305];
  assign _0527_ = sel_i[1] ? _0526_ : _0525_;
  assign _0528_ = sel_i[0] ? data_i[321] : data_i[337];
  assign _0529_ = sel_i[0] ? data_i[353] : data_i[369];
  assign _0530_ = sel_i[1] ? _0529_ : _0528_;
  assign _0531_ = sel_i[2] ? _0530_ : _0527_;
  assign _0532_ = sel_i[0] ? data_i[385] : data_i[401];
  assign _0533_ = sel_i[0] ? data_i[417] : data_i[433];
  assign _0534_ = sel_i[1] ? _0533_ : _0532_;
  assign _0535_ = sel_i[0] ? data_i[449] : data_i[465];
  assign _0536_ = sel_i[0] ? data_i[481] : data_i[497];
  assign _0537_ = sel_i[1] ? _0536_ : _0535_;
  assign _0538_ = sel_i[2] ? _0537_ : _0534_;
  assign _0539_ = sel_i[3] ? _0538_ : _0531_;
  assign data_o[17] = sel_i[4] ? _0539_ : _0524_;
  assign _0540_ = sel_i[0] ? data_i[2] : data_i[18];
  assign _0541_ = sel_i[0] ? data_i[34] : data_i[50];
  assign _0542_ = sel_i[1] ? _0541_ : _0540_;
  assign _0543_ = sel_i[0] ? data_i[66] : data_i[82];
  assign _0544_ = sel_i[0] ? data_i[98] : data_i[114];
  assign _0545_ = sel_i[1] ? _0544_ : _0543_;
  assign _0546_ = sel_i[2] ? _0545_ : _0542_;
  assign _0547_ = sel_i[0] ? data_i[130] : data_i[146];
  assign _0548_ = sel_i[0] ? data_i[162] : data_i[178];
  assign _0549_ = sel_i[1] ? _0548_ : _0547_;
  assign _0550_ = sel_i[0] ? data_i[194] : data_i[210];
  assign _0551_ = sel_i[0] ? data_i[226] : data_i[242];
  assign _0552_ = sel_i[1] ? _0551_ : _0550_;
  assign _0553_ = sel_i[2] ? _0552_ : _0549_;
  assign _0554_ = sel_i[3] ? _0553_ : _0546_;
  assign _0555_ = sel_i[0] ? data_i[258] : data_i[274];
  assign _0556_ = sel_i[0] ? data_i[290] : data_i[306];
  assign _0557_ = sel_i[1] ? _0556_ : _0555_;
  assign _0558_ = sel_i[0] ? data_i[322] : data_i[338];
  assign _0559_ = sel_i[0] ? data_i[354] : data_i[370];
  assign _0560_ = sel_i[1] ? _0559_ : _0558_;
  assign _0561_ = sel_i[2] ? _0560_ : _0557_;
  assign _0562_ = sel_i[0] ? data_i[386] : data_i[402];
  assign _0563_ = sel_i[0] ? data_i[418] : data_i[434];
  assign _0564_ = sel_i[1] ? _0563_ : _0562_;
  assign _0565_ = sel_i[0] ? data_i[450] : data_i[466];
  assign _0566_ = sel_i[0] ? data_i[482] : data_i[498];
  assign _0567_ = sel_i[1] ? _0566_ : _0565_;
  assign _0568_ = sel_i[2] ? _0567_ : _0564_;
  assign _0569_ = sel_i[3] ? _0568_ : _0561_;
  assign data_o[18] = sel_i[4] ? _0569_ : _0554_;
  assign _0570_ = sel_i[0] ? data_i[3] : data_i[19];
  assign _0571_ = sel_i[0] ? data_i[35] : data_i[51];
  assign _0572_ = sel_i[1] ? _0571_ : _0570_;
  assign _0573_ = sel_i[0] ? data_i[67] : data_i[83];
  assign _0574_ = sel_i[0] ? data_i[99] : data_i[115];
  assign _0575_ = sel_i[1] ? _0574_ : _0573_;
  assign _0576_ = sel_i[2] ? _0575_ : _0572_;
  assign _0577_ = sel_i[0] ? data_i[131] : data_i[147];
  assign _0578_ = sel_i[0] ? data_i[163] : data_i[179];
  assign _0579_ = sel_i[1] ? _0578_ : _0577_;
  assign _0580_ = sel_i[0] ? data_i[195] : data_i[211];
  assign _0581_ = sel_i[0] ? data_i[227] : data_i[243];
  assign _0582_ = sel_i[1] ? _0581_ : _0580_;
  assign _0583_ = sel_i[2] ? _0582_ : _0579_;
  assign _0584_ = sel_i[3] ? _0583_ : _0576_;
  assign _0585_ = sel_i[0] ? data_i[259] : data_i[275];
  assign _0586_ = sel_i[0] ? data_i[291] : data_i[307];
  assign _0587_ = sel_i[1] ? _0586_ : _0585_;
  assign _0588_ = sel_i[0] ? data_i[323] : data_i[339];
  assign _0589_ = sel_i[0] ? data_i[355] : data_i[371];
  assign _0590_ = sel_i[1] ? _0589_ : _0588_;
  assign _0591_ = sel_i[2] ? _0590_ : _0587_;
  assign _0592_ = sel_i[0] ? data_i[387] : data_i[403];
  assign _0593_ = sel_i[0] ? data_i[419] : data_i[435];
  assign _0594_ = sel_i[1] ? _0593_ : _0592_;
  assign _0595_ = sel_i[0] ? data_i[451] : data_i[467];
  assign _0596_ = sel_i[0] ? data_i[483] : data_i[499];
  assign _0597_ = sel_i[1] ? _0596_ : _0595_;
  assign _0598_ = sel_i[2] ? _0597_ : _0594_;
  assign _0599_ = sel_i[3] ? _0598_ : _0591_;
  assign data_o[19] = sel_i[4] ? _0599_ : _0584_;
  assign _0600_ = sel_i[0] ? data_i[4] : data_i[20];
  assign _0601_ = sel_i[0] ? data_i[36] : data_i[52];
  assign _0602_ = sel_i[1] ? _0601_ : _0600_;
  assign _0603_ = sel_i[0] ? data_i[68] : data_i[84];
  assign _0604_ = sel_i[0] ? data_i[100] : data_i[116];
  assign _0605_ = sel_i[1] ? _0604_ : _0603_;
  assign _0606_ = sel_i[2] ? _0605_ : _0602_;
  assign _0607_ = sel_i[0] ? data_i[132] : data_i[148];
  assign _0608_ = sel_i[0] ? data_i[164] : data_i[180];
  assign _0609_ = sel_i[1] ? _0608_ : _0607_;
  assign _0610_ = sel_i[0] ? data_i[196] : data_i[212];
  assign _0611_ = sel_i[0] ? data_i[228] : data_i[244];
  assign _0612_ = sel_i[1] ? _0611_ : _0610_;
  assign _0613_ = sel_i[2] ? _0612_ : _0609_;
  assign _0614_ = sel_i[3] ? _0613_ : _0606_;
  assign _0615_ = sel_i[0] ? data_i[260] : data_i[276];
  assign _0616_ = sel_i[0] ? data_i[292] : data_i[308];
  assign _0617_ = sel_i[1] ? _0616_ : _0615_;
  assign _0618_ = sel_i[0] ? data_i[324] : data_i[340];
  assign _0619_ = sel_i[0] ? data_i[356] : data_i[372];
  assign _0620_ = sel_i[1] ? _0619_ : _0618_;
  assign _0621_ = sel_i[2] ? _0620_ : _0617_;
  assign _0622_ = sel_i[0] ? data_i[388] : data_i[404];
  assign _0623_ = sel_i[0] ? data_i[420] : data_i[436];
  assign _0624_ = sel_i[1] ? _0623_ : _0622_;
  assign _0625_ = sel_i[0] ? data_i[452] : data_i[468];
  assign _0626_ = sel_i[0] ? data_i[484] : data_i[500];
  assign _0627_ = sel_i[1] ? _0626_ : _0625_;
  assign _0628_ = sel_i[2] ? _0627_ : _0624_;
  assign _0629_ = sel_i[3] ? _0628_ : _0621_;
  assign data_o[20] = sel_i[4] ? _0629_ : _0614_;
  assign _0630_ = sel_i[0] ? data_i[5] : data_i[21];
  assign _0631_ = sel_i[0] ? data_i[37] : data_i[53];
  assign _0632_ = sel_i[1] ? _0631_ : _0630_;
  assign _0633_ = sel_i[0] ? data_i[69] : data_i[85];
  assign _0634_ = sel_i[0] ? data_i[101] : data_i[117];
  assign _0635_ = sel_i[1] ? _0634_ : _0633_;
  assign _0636_ = sel_i[2] ? _0635_ : _0632_;
  assign _0637_ = sel_i[0] ? data_i[133] : data_i[149];
  assign _0638_ = sel_i[0] ? data_i[165] : data_i[181];
  assign _0639_ = sel_i[1] ? _0638_ : _0637_;
  assign _0640_ = sel_i[0] ? data_i[197] : data_i[213];
  assign _0641_ = sel_i[0] ? data_i[229] : data_i[245];
  assign _0642_ = sel_i[1] ? _0641_ : _0640_;
  assign _0643_ = sel_i[2] ? _0642_ : _0639_;
  assign _0644_ = sel_i[3] ? _0643_ : _0636_;
  assign _0645_ = sel_i[0] ? data_i[261] : data_i[277];
  assign _0646_ = sel_i[0] ? data_i[293] : data_i[309];
  assign _0647_ = sel_i[1] ? _0646_ : _0645_;
  assign _0648_ = sel_i[0] ? data_i[325] : data_i[341];
  assign _0649_ = sel_i[0] ? data_i[357] : data_i[373];
  assign _0650_ = sel_i[1] ? _0649_ : _0648_;
  assign _0651_ = sel_i[2] ? _0650_ : _0647_;
  assign _0652_ = sel_i[0] ? data_i[389] : data_i[405];
  assign _0653_ = sel_i[0] ? data_i[421] : data_i[437];
  assign _0654_ = sel_i[1] ? _0653_ : _0652_;
  assign _0655_ = sel_i[0] ? data_i[453] : data_i[469];
  assign _0656_ = sel_i[0] ? data_i[485] : data_i[501];
  assign _0657_ = sel_i[1] ? _0656_ : _0655_;
  assign _0658_ = sel_i[2] ? _0657_ : _0654_;
  assign _0659_ = sel_i[3] ? _0658_ : _0651_;
  assign data_o[21] = sel_i[4] ? _0659_ : _0644_;
  assign _0660_ = sel_i[0] ? data_i[6] : data_i[22];
  assign _0661_ = sel_i[0] ? data_i[38] : data_i[54];
  assign _0662_ = sel_i[1] ? _0661_ : _0660_;
  assign _0663_ = sel_i[0] ? data_i[70] : data_i[86];
  assign _0664_ = sel_i[0] ? data_i[102] : data_i[118];
  assign _0665_ = sel_i[1] ? _0664_ : _0663_;
  assign _0666_ = sel_i[2] ? _0665_ : _0662_;
  assign _0667_ = sel_i[0] ? data_i[134] : data_i[150];
  assign _0668_ = sel_i[0] ? data_i[166] : data_i[182];
  assign _0669_ = sel_i[1] ? _0668_ : _0667_;
  assign _0670_ = sel_i[0] ? data_i[198] : data_i[214];
  assign _0671_ = sel_i[0] ? data_i[230] : data_i[246];
  assign _0672_ = sel_i[1] ? _0671_ : _0670_;
  assign _0673_ = sel_i[2] ? _0672_ : _0669_;
  assign _0674_ = sel_i[3] ? _0673_ : _0666_;
  assign _0675_ = sel_i[0] ? data_i[262] : data_i[278];
  assign _0676_ = sel_i[0] ? data_i[294] : data_i[310];
  assign _0677_ = sel_i[1] ? _0676_ : _0675_;
  assign _0678_ = sel_i[0] ? data_i[326] : data_i[342];
  assign _0679_ = sel_i[0] ? data_i[358] : data_i[374];
  assign _0680_ = sel_i[1] ? _0679_ : _0678_;
  assign _0681_ = sel_i[2] ? _0680_ : _0677_;
  assign _0682_ = sel_i[0] ? data_i[390] : data_i[406];
  assign _0683_ = sel_i[0] ? data_i[422] : data_i[438];
  assign _0684_ = sel_i[1] ? _0683_ : _0682_;
  assign _0685_ = sel_i[0] ? data_i[454] : data_i[470];
  assign _0686_ = sel_i[0] ? data_i[486] : data_i[502];
  assign _0687_ = sel_i[1] ? _0686_ : _0685_;
  assign _0688_ = sel_i[2] ? _0687_ : _0684_;
  assign _0689_ = sel_i[3] ? _0688_ : _0681_;
  assign data_o[22] = sel_i[4] ? _0689_ : _0674_;
  assign _0690_ = sel_i[0] ? data_i[7] : data_i[23];
  assign _0691_ = sel_i[0] ? data_i[39] : data_i[55];
  assign _0692_ = sel_i[1] ? _0691_ : _0690_;
  assign _0693_ = sel_i[0] ? data_i[71] : data_i[87];
  assign _0694_ = sel_i[0] ? data_i[103] : data_i[119];
  assign _0695_ = sel_i[1] ? _0694_ : _0693_;
  assign _0696_ = sel_i[2] ? _0695_ : _0692_;
  assign _0697_ = sel_i[0] ? data_i[135] : data_i[151];
  assign _0698_ = sel_i[0] ? data_i[167] : data_i[183];
  assign _0699_ = sel_i[1] ? _0698_ : _0697_;
  assign _0700_ = sel_i[0] ? data_i[199] : data_i[215];
  assign _0701_ = sel_i[0] ? data_i[231] : data_i[247];
  assign _0702_ = sel_i[1] ? _0701_ : _0700_;
  assign _0703_ = sel_i[2] ? _0702_ : _0699_;
  assign _0704_ = sel_i[3] ? _0703_ : _0696_;
  assign _0705_ = sel_i[0] ? data_i[263] : data_i[279];
  assign _0706_ = sel_i[0] ? data_i[295] : data_i[311];
  assign _0707_ = sel_i[1] ? _0706_ : _0705_;
  assign _0708_ = sel_i[0] ? data_i[327] : data_i[343];
  assign _0709_ = sel_i[0] ? data_i[359] : data_i[375];
  assign _0710_ = sel_i[1] ? _0709_ : _0708_;
  assign _0711_ = sel_i[2] ? _0710_ : _0707_;
  assign _0712_ = sel_i[0] ? data_i[391] : data_i[407];
  assign _0713_ = sel_i[0] ? data_i[423] : data_i[439];
  assign _0714_ = sel_i[1] ? _0713_ : _0712_;
  assign _0715_ = sel_i[0] ? data_i[455] : data_i[471];
  assign _0716_ = sel_i[0] ? data_i[487] : data_i[503];
  assign _0717_ = sel_i[1] ? _0716_ : _0715_;
  assign _0718_ = sel_i[2] ? _0717_ : _0714_;
  assign _0719_ = sel_i[3] ? _0718_ : _0711_;
  assign data_o[23] = sel_i[4] ? _0719_ : _0704_;
  assign _0720_ = sel_i[0] ? data_i[8] : data_i[24];
  assign _0721_ = sel_i[0] ? data_i[40] : data_i[56];
  assign _0722_ = sel_i[1] ? _0721_ : _0720_;
  assign _0723_ = sel_i[0] ? data_i[72] : data_i[88];
  assign _0724_ = sel_i[0] ? data_i[104] : data_i[120];
  assign _0725_ = sel_i[1] ? _0724_ : _0723_;
  assign _0726_ = sel_i[2] ? _0725_ : _0722_;
  assign _0727_ = sel_i[0] ? data_i[136] : data_i[152];
  assign _0728_ = sel_i[0] ? data_i[168] : data_i[184];
  assign _0729_ = sel_i[1] ? _0728_ : _0727_;
  assign _0730_ = sel_i[0] ? data_i[200] : data_i[216];
  assign _0731_ = sel_i[0] ? data_i[232] : data_i[248];
  assign _0732_ = sel_i[1] ? _0731_ : _0730_;
  assign _0733_ = sel_i[2] ? _0732_ : _0729_;
  assign _0734_ = sel_i[3] ? _0733_ : _0726_;
  assign _0735_ = sel_i[0] ? data_i[264] : data_i[280];
  assign _0736_ = sel_i[0] ? data_i[296] : data_i[312];
  assign _0737_ = sel_i[1] ? _0736_ : _0735_;
  assign _0738_ = sel_i[0] ? data_i[328] : data_i[344];
  assign _0739_ = sel_i[0] ? data_i[360] : data_i[376];
  assign _0740_ = sel_i[1] ? _0739_ : _0738_;
  assign _0741_ = sel_i[2] ? _0740_ : _0737_;
  assign _0742_ = sel_i[0] ? data_i[392] : data_i[408];
  assign _0743_ = sel_i[0] ? data_i[424] : data_i[440];
  assign _0744_ = sel_i[1] ? _0743_ : _0742_;
  assign _0745_ = sel_i[0] ? data_i[456] : data_i[472];
  assign _0746_ = sel_i[0] ? data_i[488] : data_i[504];
  assign _0747_ = sel_i[1] ? _0746_ : _0745_;
  assign _0748_ = sel_i[2] ? _0747_ : _0744_;
  assign _0749_ = sel_i[3] ? _0748_ : _0741_;
  assign data_o[24] = sel_i[4] ? _0749_ : _0734_;
  assign _0750_ = sel_i[0] ? data_i[9] : data_i[25];
  assign _0751_ = sel_i[0] ? data_i[41] : data_i[57];
  assign _0752_ = sel_i[1] ? _0751_ : _0750_;
  assign _0753_ = sel_i[0] ? data_i[73] : data_i[89];
  assign _0754_ = sel_i[0] ? data_i[105] : data_i[121];
  assign _0755_ = sel_i[1] ? _0754_ : _0753_;
  assign _0756_ = sel_i[2] ? _0755_ : _0752_;
  assign _0757_ = sel_i[0] ? data_i[137] : data_i[153];
  assign _0758_ = sel_i[0] ? data_i[169] : data_i[185];
  assign _0759_ = sel_i[1] ? _0758_ : _0757_;
  assign _0760_ = sel_i[0] ? data_i[201] : data_i[217];
  assign _0761_ = sel_i[0] ? data_i[233] : data_i[249];
  assign _0762_ = sel_i[1] ? _0761_ : _0760_;
  assign _0763_ = sel_i[2] ? _0762_ : _0759_;
  assign _0764_ = sel_i[3] ? _0763_ : _0756_;
  assign _0765_ = sel_i[0] ? data_i[265] : data_i[281];
  assign _0766_ = sel_i[0] ? data_i[297] : data_i[313];
  assign _0767_ = sel_i[1] ? _0766_ : _0765_;
  assign _0768_ = sel_i[0] ? data_i[329] : data_i[345];
  assign _0769_ = sel_i[0] ? data_i[361] : data_i[377];
  assign _0770_ = sel_i[1] ? _0769_ : _0768_;
  assign _0771_ = sel_i[2] ? _0770_ : _0767_;
  assign _0772_ = sel_i[0] ? data_i[393] : data_i[409];
  assign _0773_ = sel_i[0] ? data_i[425] : data_i[441];
  assign _0774_ = sel_i[1] ? _0773_ : _0772_;
  assign _0775_ = sel_i[0] ? data_i[457] : data_i[473];
  assign _0776_ = sel_i[0] ? data_i[489] : data_i[505];
  assign _0777_ = sel_i[1] ? _0776_ : _0775_;
  assign _0778_ = sel_i[2] ? _0777_ : _0774_;
  assign _0779_ = sel_i[3] ? _0778_ : _0771_;
  assign data_o[25] = sel_i[4] ? _0779_ : _0764_;
  assign _0780_ = sel_i[0] ? data_i[10] : data_i[26];
  assign _0781_ = sel_i[0] ? data_i[42] : data_i[58];
  assign _0782_ = sel_i[1] ? _0781_ : _0780_;
  assign _0783_ = sel_i[0] ? data_i[74] : data_i[90];
  assign _0784_ = sel_i[0] ? data_i[106] : data_i[122];
  assign _0785_ = sel_i[1] ? _0784_ : _0783_;
  assign _0786_ = sel_i[2] ? _0785_ : _0782_;
  assign _0787_ = sel_i[0] ? data_i[138] : data_i[154];
  assign _0788_ = sel_i[0] ? data_i[170] : data_i[186];
  assign _0789_ = sel_i[1] ? _0788_ : _0787_;
  assign _0790_ = sel_i[0] ? data_i[202] : data_i[218];
  assign _0791_ = sel_i[0] ? data_i[234] : data_i[250];
  assign _0792_ = sel_i[1] ? _0791_ : _0790_;
  assign _0793_ = sel_i[2] ? _0792_ : _0789_;
  assign _0794_ = sel_i[3] ? _0793_ : _0786_;
  assign _0795_ = sel_i[0] ? data_i[266] : data_i[282];
  assign _0796_ = sel_i[0] ? data_i[298] : data_i[314];
  assign _0797_ = sel_i[1] ? _0796_ : _0795_;
  assign _0798_ = sel_i[0] ? data_i[330] : data_i[346];
  assign _0799_ = sel_i[0] ? data_i[362] : data_i[378];
  assign _0800_ = sel_i[1] ? _0799_ : _0798_;
  assign _0801_ = sel_i[2] ? _0800_ : _0797_;
  assign _0802_ = sel_i[0] ? data_i[394] : data_i[410];
  assign _0803_ = sel_i[0] ? data_i[426] : data_i[442];
  assign _0804_ = sel_i[1] ? _0803_ : _0802_;
  assign _0805_ = sel_i[0] ? data_i[458] : data_i[474];
  assign _0806_ = sel_i[0] ? data_i[490] : data_i[506];
  assign _0807_ = sel_i[1] ? _0806_ : _0805_;
  assign _0808_ = sel_i[2] ? _0807_ : _0804_;
  assign _0809_ = sel_i[3] ? _0808_ : _0801_;
  assign data_o[26] = sel_i[4] ? _0809_ : _0794_;
  assign _0810_ = sel_i[0] ? data_i[11] : data_i[27];
  assign _0811_ = sel_i[0] ? data_i[43] : data_i[59];
  assign _0812_ = sel_i[1] ? _0811_ : _0810_;
  assign _0813_ = sel_i[0] ? data_i[75] : data_i[91];
  assign _0814_ = sel_i[0] ? data_i[107] : data_i[123];
  assign _0815_ = sel_i[1] ? _0814_ : _0813_;
  assign _0816_ = sel_i[2] ? _0815_ : _0812_;
  assign _0817_ = sel_i[0] ? data_i[139] : data_i[155];
  assign _0818_ = sel_i[0] ? data_i[171] : data_i[187];
  assign _0819_ = sel_i[1] ? _0818_ : _0817_;
  assign _0820_ = sel_i[0] ? data_i[203] : data_i[219];
  assign _0821_ = sel_i[0] ? data_i[235] : data_i[251];
  assign _0822_ = sel_i[1] ? _0821_ : _0820_;
  assign _0823_ = sel_i[2] ? _0822_ : _0819_;
  assign _0824_ = sel_i[3] ? _0823_ : _0816_;
  assign _0825_ = sel_i[0] ? data_i[267] : data_i[283];
  assign _0826_ = sel_i[0] ? data_i[299] : data_i[315];
  assign _0827_ = sel_i[1] ? _0826_ : _0825_;
  assign _0828_ = sel_i[0] ? data_i[331] : data_i[347];
  assign _0829_ = sel_i[0] ? data_i[363] : data_i[379];
  assign _0830_ = sel_i[1] ? _0829_ : _0828_;
  assign _0831_ = sel_i[2] ? _0830_ : _0827_;
  assign _0832_ = sel_i[0] ? data_i[395] : data_i[411];
  assign _0833_ = sel_i[0] ? data_i[427] : data_i[443];
  assign _0834_ = sel_i[1] ? _0833_ : _0832_;
  assign _0835_ = sel_i[0] ? data_i[459] : data_i[475];
  assign _0836_ = sel_i[0] ? data_i[491] : data_i[507];
  assign _0837_ = sel_i[1] ? _0836_ : _0835_;
  assign _0838_ = sel_i[2] ? _0837_ : _0834_;
  assign _0839_ = sel_i[3] ? _0838_ : _0831_;
  assign data_o[27] = sel_i[4] ? _0839_ : _0824_;
  assign _0840_ = sel_i[0] ? data_i[12] : data_i[28];
  assign _0841_ = sel_i[0] ? data_i[44] : data_i[60];
  assign _0842_ = sel_i[1] ? _0841_ : _0840_;
  assign _0843_ = sel_i[0] ? data_i[76] : data_i[92];
  assign _0844_ = sel_i[0] ? data_i[108] : data_i[124];
  assign _0845_ = sel_i[1] ? _0844_ : _0843_;
  assign _0846_ = sel_i[2] ? _0845_ : _0842_;
  assign _0847_ = sel_i[0] ? data_i[140] : data_i[156];
  assign _0848_ = sel_i[0] ? data_i[172] : data_i[188];
  assign _0849_ = sel_i[1] ? _0848_ : _0847_;
  assign _0850_ = sel_i[0] ? data_i[204] : data_i[220];
  assign _0851_ = sel_i[0] ? data_i[236] : data_i[252];
  assign _0852_ = sel_i[1] ? _0851_ : _0850_;
  assign _0853_ = sel_i[2] ? _0852_ : _0849_;
  assign _0854_ = sel_i[3] ? _0853_ : _0846_;
  assign _0855_ = sel_i[0] ? data_i[268] : data_i[284];
  assign _0856_ = sel_i[0] ? data_i[300] : data_i[316];
  assign _0857_ = sel_i[1] ? _0856_ : _0855_;
  assign _0858_ = sel_i[0] ? data_i[332] : data_i[348];
  assign _0859_ = sel_i[0] ? data_i[364] : data_i[380];
  assign _0860_ = sel_i[1] ? _0859_ : _0858_;
  assign _0861_ = sel_i[2] ? _0860_ : _0857_;
  assign _0862_ = sel_i[0] ? data_i[396] : data_i[412];
  assign _0863_ = sel_i[0] ? data_i[428] : data_i[444];
  assign _0864_ = sel_i[1] ? _0863_ : _0862_;
  assign _0865_ = sel_i[0] ? data_i[460] : data_i[476];
  assign _0866_ = sel_i[0] ? data_i[492] : data_i[508];
  assign _0867_ = sel_i[1] ? _0866_ : _0865_;
  assign _0868_ = sel_i[2] ? _0867_ : _0864_;
  assign _0869_ = sel_i[3] ? _0868_ : _0861_;
  assign data_o[28] = sel_i[4] ? _0869_ : _0854_;
  assign _0870_ = sel_i[0] ? data_i[13] : data_i[29];
  assign _0871_ = sel_i[0] ? data_i[45] : data_i[61];
  assign _0872_ = sel_i[1] ? _0871_ : _0870_;
  assign _0873_ = sel_i[0] ? data_i[77] : data_i[93];
  assign _0874_ = sel_i[0] ? data_i[109] : data_i[125];
  assign _0875_ = sel_i[1] ? _0874_ : _0873_;
  assign _0876_ = sel_i[2] ? _0875_ : _0872_;
  assign _0877_ = sel_i[0] ? data_i[141] : data_i[157];
  assign _0878_ = sel_i[0] ? data_i[173] : data_i[189];
  assign _0879_ = sel_i[1] ? _0878_ : _0877_;
  assign _0880_ = sel_i[0] ? data_i[205] : data_i[221];
  assign _0881_ = sel_i[0] ? data_i[237] : data_i[253];
  assign _0882_ = sel_i[1] ? _0881_ : _0880_;
  assign _0883_ = sel_i[2] ? _0882_ : _0879_;
  assign _0884_ = sel_i[3] ? _0883_ : _0876_;
  assign _0885_ = sel_i[0] ? data_i[269] : data_i[285];
  assign _0886_ = sel_i[0] ? data_i[301] : data_i[317];
  assign _0887_ = sel_i[1] ? _0886_ : _0885_;
  assign _0888_ = sel_i[0] ? data_i[333] : data_i[349];
  assign _0889_ = sel_i[0] ? data_i[365] : data_i[381];
  assign _0890_ = sel_i[1] ? _0889_ : _0888_;
  assign _0891_ = sel_i[2] ? _0890_ : _0887_;
  assign _0892_ = sel_i[0] ? data_i[397] : data_i[413];
  assign _0893_ = sel_i[0] ? data_i[429] : data_i[445];
  assign _0894_ = sel_i[1] ? _0893_ : _0892_;
  assign _0895_ = sel_i[0] ? data_i[461] : data_i[477];
  assign _0896_ = sel_i[0] ? data_i[493] : data_i[509];
  assign _0897_ = sel_i[1] ? _0896_ : _0895_;
  assign _0898_ = sel_i[2] ? _0897_ : _0894_;
  assign _0899_ = sel_i[3] ? _0898_ : _0891_;
  assign data_o[29] = sel_i[4] ? _0899_ : _0884_;
  assign _0900_ = sel_i[0] ? data_i[14] : data_i[30];
  assign _0901_ = sel_i[0] ? data_i[46] : data_i[62];
  assign _0902_ = sel_i[1] ? _0901_ : _0900_;
  assign _0903_ = sel_i[0] ? data_i[78] : data_i[94];
  assign _0904_ = sel_i[0] ? data_i[110] : data_i[126];
  assign _0905_ = sel_i[1] ? _0904_ : _0903_;
  assign _0906_ = sel_i[2] ? _0905_ : _0902_;
  assign _0907_ = sel_i[0] ? data_i[142] : data_i[158];
  assign _0908_ = sel_i[0] ? data_i[174] : data_i[190];
  assign _0909_ = sel_i[1] ? _0908_ : _0907_;
  assign _0910_ = sel_i[0] ? data_i[206] : data_i[222];
  assign _0911_ = sel_i[0] ? data_i[238] : data_i[254];
  assign _0912_ = sel_i[1] ? _0911_ : _0910_;
  assign _0913_ = sel_i[2] ? _0912_ : _0909_;
  assign _0914_ = sel_i[3] ? _0913_ : _0906_;
  assign _0915_ = sel_i[0] ? data_i[270] : data_i[286];
  assign _0916_ = sel_i[0] ? data_i[302] : data_i[318];
  assign _0917_ = sel_i[1] ? _0916_ : _0915_;
  assign _0918_ = sel_i[0] ? data_i[334] : data_i[350];
  assign _0919_ = sel_i[0] ? data_i[366] : data_i[382];
  assign _0920_ = sel_i[1] ? _0919_ : _0918_;
  assign _0921_ = sel_i[2] ? _0920_ : _0917_;
  assign _0922_ = sel_i[0] ? data_i[398] : data_i[414];
  assign _0923_ = sel_i[0] ? data_i[430] : data_i[446];
  assign _0924_ = sel_i[1] ? _0923_ : _0922_;
  assign _0925_ = sel_i[0] ? data_i[462] : data_i[478];
  assign _0926_ = sel_i[0] ? data_i[494] : data_i[510];
  assign _0927_ = sel_i[1] ? _0926_ : _0925_;
  assign _0928_ = sel_i[2] ? _0927_ : _0924_;
  assign _0929_ = sel_i[3] ? _0928_ : _0921_;
  assign data_o[30] = sel_i[4] ? _0929_ : _0914_;
  assign _0930_ = sel_i[0] ? data_i[15] : data_i[31];
  assign _0931_ = sel_i[0] ? data_i[47] : data_i[63];
  assign _0932_ = sel_i[1] ? _0931_ : _0930_;
  assign _0933_ = sel_i[0] ? data_i[79] : data_i[95];
  assign _0934_ = sel_i[0] ? data_i[111] : data_i[127];
  assign _0935_ = sel_i[1] ? _0934_ : _0933_;
  assign _0936_ = sel_i[2] ? _0935_ : _0932_;
  assign _0937_ = sel_i[0] ? data_i[143] : data_i[159];
  assign _0938_ = sel_i[0] ? data_i[175] : data_i[191];
  assign _0939_ = sel_i[1] ? _0938_ : _0937_;
  assign _0940_ = sel_i[0] ? data_i[207] : data_i[223];
  assign _0941_ = sel_i[0] ? data_i[239] : data_i[255];
  assign _0942_ = sel_i[1] ? _0941_ : _0940_;
  assign _0943_ = sel_i[2] ? _0942_ : _0939_;
  assign _0944_ = sel_i[3] ? _0943_ : _0936_;
  assign _0945_ = sel_i[0] ? data_i[271] : data_i[287];
  assign _0946_ = sel_i[0] ? data_i[303] : data_i[319];
  assign _0947_ = sel_i[1] ? _0946_ : _0945_;
  assign _0948_ = sel_i[0] ? data_i[335] : data_i[351];
  assign _0949_ = sel_i[0] ? data_i[367] : data_i[383];
  assign _0950_ = sel_i[1] ? _0949_ : _0948_;
  assign _0951_ = sel_i[2] ? _0950_ : _0947_;
  assign _0952_ = sel_i[0] ? data_i[399] : data_i[415];
  assign _0953_ = sel_i[0] ? data_i[431] : data_i[447];
  assign _0954_ = sel_i[1] ? _0953_ : _0952_;
  assign _0955_ = sel_i[0] ? data_i[463] : data_i[479];
  assign _0956_ = sel_i[0] ? data_i[495] : data_i[511];
  assign _0957_ = sel_i[1] ? _0956_ : _0955_;
  assign _0958_ = sel_i[2] ? _0957_ : _0954_;
  assign _0959_ = sel_i[3] ? _0958_ : _0951_;
  assign data_o[31] = sel_i[4] ? _0959_ : _0944_;
  assign _0960_ = sel_i[1] ? _0000_ : _0001_;
  assign _0961_ = sel_i[1] ? _0003_ : _0004_;
  assign _0962_ = sel_i[2] ? _0961_ : _0960_;
  assign _0963_ = sel_i[1] ? _0007_ : _0008_;
  assign _0964_ = sel_i[1] ? _0010_ : _0011_;
  assign _0965_ = sel_i[2] ? _0964_ : _0963_;
  assign _0966_ = sel_i[3] ? _0965_ : _0962_;
  assign _0967_ = sel_i[1] ? _0015_ : _0016_;
  assign _0968_ = sel_i[1] ? _0018_ : _0019_;
  assign _0969_ = sel_i[2] ? _0968_ : _0967_;
  assign _0970_ = sel_i[1] ? _0022_ : _0023_;
  assign _0971_ = sel_i[1] ? _0025_ : _0026_;
  assign _0972_ = sel_i[2] ? _0971_ : _0970_;
  assign _0973_ = sel_i[3] ? _0972_ : _0969_;
  assign data_o[32] = sel_i[4] ? _0973_ : _0966_;
  assign _0974_ = sel_i[1] ? _0030_ : _0031_;
  assign _0975_ = sel_i[1] ? _0033_ : _0034_;
  assign _0976_ = sel_i[2] ? _0975_ : _0974_;
  assign _0977_ = sel_i[1] ? _0037_ : _0038_;
  assign _0978_ = sel_i[1] ? _0040_ : _0041_;
  assign _0979_ = sel_i[2] ? _0978_ : _0977_;
  assign _0980_ = sel_i[3] ? _0979_ : _0976_;
  assign _0981_ = sel_i[1] ? _0045_ : _0046_;
  assign _0982_ = sel_i[1] ? _0048_ : _0049_;
  assign _0983_ = sel_i[2] ? _0982_ : _0981_;
  assign _0984_ = sel_i[1] ? _0052_ : _0053_;
  assign _0985_ = sel_i[1] ? _0055_ : _0056_;
  assign _0986_ = sel_i[2] ? _0985_ : _0984_;
  assign _0987_ = sel_i[3] ? _0986_ : _0983_;
  assign data_o[33] = sel_i[4] ? _0987_ : _0980_;
  assign _0988_ = sel_i[1] ? _0060_ : _0061_;
  assign _0989_ = sel_i[1] ? _0063_ : _0064_;
  assign _0990_ = sel_i[2] ? _0989_ : _0988_;
  assign _0991_ = sel_i[1] ? _0067_ : _0068_;
  assign _0992_ = sel_i[1] ? _0070_ : _0071_;
  assign _0993_ = sel_i[2] ? _0992_ : _0991_;
  assign _0994_ = sel_i[3] ? _0993_ : _0990_;
  assign _0995_ = sel_i[1] ? _0075_ : _0076_;
  assign _0996_ = sel_i[1] ? _0078_ : _0079_;
  assign _0997_ = sel_i[2] ? _0996_ : _0995_;
  assign _0998_ = sel_i[1] ? _0082_ : _0083_;
  assign _0999_ = sel_i[1] ? _0085_ : _0086_;
  assign _1000_ = sel_i[2] ? _0999_ : _0998_;
  assign _1001_ = sel_i[3] ? _1000_ : _0997_;
  assign data_o[34] = sel_i[4] ? _1001_ : _0994_;
  assign _1002_ = sel_i[1] ? _0090_ : _0091_;
  assign _1003_ = sel_i[1] ? _0093_ : _0094_;
  assign _1004_ = sel_i[2] ? _1003_ : _1002_;
  assign _1005_ = sel_i[1] ? _0097_ : _0098_;
  assign _1006_ = sel_i[1] ? _0100_ : _0101_;
  assign _1007_ = sel_i[2] ? _1006_ : _1005_;
  assign _1008_ = sel_i[3] ? _1007_ : _1004_;
  assign _1009_ = sel_i[1] ? _0105_ : _0106_;
  assign _1010_ = sel_i[1] ? _0108_ : _0109_;
  assign _1011_ = sel_i[2] ? _1010_ : _1009_;
  assign _1012_ = sel_i[1] ? _0112_ : _0113_;
  assign _1013_ = sel_i[1] ? _0115_ : _0116_;
  assign _1014_ = sel_i[2] ? _1013_ : _1012_;
  assign _1015_ = sel_i[3] ? _1014_ : _1011_;
  assign data_o[35] = sel_i[4] ? _1015_ : _1008_;
  assign _1016_ = sel_i[1] ? _0120_ : _0121_;
  assign _1017_ = sel_i[1] ? _0123_ : _0124_;
  assign _1018_ = sel_i[2] ? _1017_ : _1016_;
  assign _1019_ = sel_i[1] ? _0127_ : _0128_;
  assign _1020_ = sel_i[1] ? _0130_ : _0131_;
  assign _1021_ = sel_i[2] ? _1020_ : _1019_;
  assign _1022_ = sel_i[3] ? _1021_ : _1018_;
  assign _1023_ = sel_i[1] ? _0135_ : _0136_;
  assign _1024_ = sel_i[1] ? _0138_ : _0139_;
  assign _1025_ = sel_i[2] ? _1024_ : _1023_;
  assign _1026_ = sel_i[1] ? _0142_ : _0143_;
  assign _1027_ = sel_i[1] ? _0145_ : _0146_;
  assign _1028_ = sel_i[2] ? _1027_ : _1026_;
  assign _1029_ = sel_i[3] ? _1028_ : _1025_;
  assign data_o[36] = sel_i[4] ? _1029_ : _1022_;
  assign _1030_ = sel_i[1] ? _0150_ : _0151_;
  assign _1031_ = sel_i[1] ? _0153_ : _0154_;
  assign _1032_ = sel_i[2] ? _1031_ : _1030_;
  assign _1033_ = sel_i[1] ? _0157_ : _0158_;
  assign _1034_ = sel_i[1] ? _0160_ : _0161_;
  assign _1035_ = sel_i[2] ? _1034_ : _1033_;
  assign _1036_ = sel_i[3] ? _1035_ : _1032_;
  assign _1037_ = sel_i[1] ? _0165_ : _0166_;
  assign _1038_ = sel_i[1] ? _0168_ : _0169_;
  assign _1039_ = sel_i[2] ? _1038_ : _1037_;
  assign _1040_ = sel_i[1] ? _0172_ : _0173_;
  assign _1041_ = sel_i[1] ? _0175_ : _0176_;
  assign _1042_ = sel_i[2] ? _1041_ : _1040_;
  assign _1043_ = sel_i[3] ? _1042_ : _1039_;
  assign data_o[37] = sel_i[4] ? _1043_ : _1036_;
  assign _1044_ = sel_i[1] ? _0180_ : _0181_;
  assign _1045_ = sel_i[1] ? _0183_ : _0184_;
  assign _1046_ = sel_i[2] ? _1045_ : _1044_;
  assign _1047_ = sel_i[1] ? _0187_ : _0188_;
  assign _1048_ = sel_i[1] ? _0190_ : _0191_;
  assign _1049_ = sel_i[2] ? _1048_ : _1047_;
  assign _1050_ = sel_i[3] ? _1049_ : _1046_;
  assign _1051_ = sel_i[1] ? _0195_ : _0196_;
  assign _1052_ = sel_i[1] ? _0198_ : _0199_;
  assign _1053_ = sel_i[2] ? _1052_ : _1051_;
  assign _1054_ = sel_i[1] ? _0202_ : _0203_;
  assign _1055_ = sel_i[1] ? _0205_ : _0206_;
  assign _1056_ = sel_i[2] ? _1055_ : _1054_;
  assign _1057_ = sel_i[3] ? _1056_ : _1053_;
  assign data_o[38] = sel_i[4] ? _1057_ : _1050_;
  assign _1058_ = sel_i[1] ? _0210_ : _0211_;
  assign _1059_ = sel_i[1] ? _0213_ : _0214_;
  assign _1060_ = sel_i[2] ? _1059_ : _1058_;
  assign _1061_ = sel_i[1] ? _0217_ : _0218_;
  assign _1062_ = sel_i[1] ? _0220_ : _0221_;
  assign _1063_ = sel_i[2] ? _1062_ : _1061_;
  assign _1064_ = sel_i[3] ? _1063_ : _1060_;
  assign _1065_ = sel_i[1] ? _0225_ : _0226_;
  assign _1066_ = sel_i[1] ? _0228_ : _0229_;
  assign _1067_ = sel_i[2] ? _1066_ : _1065_;
  assign _1068_ = sel_i[1] ? _0232_ : _0233_;
  assign _1069_ = sel_i[1] ? _0235_ : _0236_;
  assign _1070_ = sel_i[2] ? _1069_ : _1068_;
  assign _1071_ = sel_i[3] ? _1070_ : _1067_;
  assign data_o[39] = sel_i[4] ? _1071_ : _1064_;
  assign _1072_ = sel_i[1] ? _0240_ : _0241_;
  assign _1073_ = sel_i[1] ? _0243_ : _0244_;
  assign _1074_ = sel_i[2] ? _1073_ : _1072_;
  assign _1075_ = sel_i[1] ? _0247_ : _0248_;
  assign _1076_ = sel_i[1] ? _0250_ : _0251_;
  assign _1077_ = sel_i[2] ? _1076_ : _1075_;
  assign _1078_ = sel_i[3] ? _1077_ : _1074_;
  assign _1079_ = sel_i[1] ? _0255_ : _0256_;
  assign _1080_ = sel_i[1] ? _0258_ : _0259_;
  assign _1081_ = sel_i[2] ? _1080_ : _1079_;
  assign _1082_ = sel_i[1] ? _0262_ : _0263_;
  assign _1083_ = sel_i[1] ? _0265_ : _0266_;
  assign _1084_ = sel_i[2] ? _1083_ : _1082_;
  assign _1085_ = sel_i[3] ? _1084_ : _1081_;
  assign data_o[40] = sel_i[4] ? _1085_ : _1078_;
  assign _1086_ = sel_i[1] ? _0270_ : _0271_;
  assign _1087_ = sel_i[1] ? _0273_ : _0274_;
  assign _1088_ = sel_i[2] ? _1087_ : _1086_;
  assign _1089_ = sel_i[1] ? _0277_ : _0278_;
  assign _1090_ = sel_i[1] ? _0280_ : _0281_;
  assign _1091_ = sel_i[2] ? _1090_ : _1089_;
  assign _1092_ = sel_i[3] ? _1091_ : _1088_;
  assign _1093_ = sel_i[1] ? _0285_ : _0286_;
  assign _1094_ = sel_i[1] ? _0288_ : _0289_;
  assign _1095_ = sel_i[2] ? _1094_ : _1093_;
  assign _1096_ = sel_i[1] ? _0292_ : _0293_;
  assign _1097_ = sel_i[1] ? _0295_ : _0296_;
  assign _1098_ = sel_i[2] ? _1097_ : _1096_;
  assign _1099_ = sel_i[3] ? _1098_ : _1095_;
  assign data_o[41] = sel_i[4] ? _1099_ : _1092_;
  assign _1100_ = sel_i[1] ? _0300_ : _0301_;
  assign _1101_ = sel_i[1] ? _0303_ : _0304_;
  assign _1102_ = sel_i[2] ? _1101_ : _1100_;
  assign _1103_ = sel_i[1] ? _0307_ : _0308_;
  assign _1104_ = sel_i[1] ? _0310_ : _0311_;
  assign _1105_ = sel_i[2] ? _1104_ : _1103_;
  assign _1106_ = sel_i[3] ? _1105_ : _1102_;
  assign _1107_ = sel_i[1] ? _0315_ : _0316_;
  assign _1108_ = sel_i[1] ? _0318_ : _0319_;
  assign _1109_ = sel_i[2] ? _1108_ : _1107_;
  assign _1110_ = sel_i[1] ? _0322_ : _0323_;
  assign _1111_ = sel_i[1] ? _0325_ : _0326_;
  assign _1112_ = sel_i[2] ? _1111_ : _1110_;
  assign _1113_ = sel_i[3] ? _1112_ : _1109_;
  assign data_o[42] = sel_i[4] ? _1113_ : _1106_;
  assign _1114_ = sel_i[1] ? _0330_ : _0331_;
  assign _1115_ = sel_i[1] ? _0333_ : _0334_;
  assign _1116_ = sel_i[2] ? _1115_ : _1114_;
  assign _1117_ = sel_i[1] ? _0337_ : _0338_;
  assign _1118_ = sel_i[1] ? _0340_ : _0341_;
  assign _1119_ = sel_i[2] ? _1118_ : _1117_;
  assign _1120_ = sel_i[3] ? _1119_ : _1116_;
  assign _1121_ = sel_i[1] ? _0345_ : _0346_;
  assign _1122_ = sel_i[1] ? _0348_ : _0349_;
  assign _1123_ = sel_i[2] ? _1122_ : _1121_;
  assign _1124_ = sel_i[1] ? _0352_ : _0353_;
  assign _1125_ = sel_i[1] ? _0355_ : _0356_;
  assign _1126_ = sel_i[2] ? _1125_ : _1124_;
  assign _1127_ = sel_i[3] ? _1126_ : _1123_;
  assign data_o[43] = sel_i[4] ? _1127_ : _1120_;
  assign _1128_ = sel_i[1] ? _0360_ : _0361_;
  assign _1129_ = sel_i[1] ? _0363_ : _0364_;
  assign _1130_ = sel_i[2] ? _1129_ : _1128_;
  assign _1131_ = sel_i[1] ? _0367_ : _0368_;
  assign _1132_ = sel_i[1] ? _0370_ : _0371_;
  assign _1133_ = sel_i[2] ? _1132_ : _1131_;
  assign _1134_ = sel_i[3] ? _1133_ : _1130_;
  assign _1135_ = sel_i[1] ? _0375_ : _0376_;
  assign _1136_ = sel_i[1] ? _0378_ : _0379_;
  assign _1137_ = sel_i[2] ? _1136_ : _1135_;
  assign _1138_ = sel_i[1] ? _0382_ : _0383_;
  assign _1139_ = sel_i[1] ? _0385_ : _0386_;
  assign _1140_ = sel_i[2] ? _1139_ : _1138_;
  assign _1141_ = sel_i[3] ? _1140_ : _1137_;
  assign data_o[44] = sel_i[4] ? _1141_ : _1134_;
  assign _1142_ = sel_i[1] ? _0390_ : _0391_;
  assign _1143_ = sel_i[1] ? _0393_ : _0394_;
  assign _1144_ = sel_i[2] ? _1143_ : _1142_;
  assign _1145_ = sel_i[1] ? _0397_ : _0398_;
  assign _1146_ = sel_i[1] ? _0400_ : _0401_;
  assign _1147_ = sel_i[2] ? _1146_ : _1145_;
  assign _1148_ = sel_i[3] ? _1147_ : _1144_;
  assign _1149_ = sel_i[1] ? _0405_ : _0406_;
  assign _1150_ = sel_i[1] ? _0408_ : _0409_;
  assign _1151_ = sel_i[2] ? _1150_ : _1149_;
  assign _1152_ = sel_i[1] ? _0412_ : _0413_;
  assign _1153_ = sel_i[1] ? _0415_ : _0416_;
  assign _1154_ = sel_i[2] ? _1153_ : _1152_;
  assign _1155_ = sel_i[3] ? _1154_ : _1151_;
  assign data_o[45] = sel_i[4] ? _1155_ : _1148_;
  assign _1156_ = sel_i[1] ? _0420_ : _0421_;
  assign _1157_ = sel_i[1] ? _0423_ : _0424_;
  assign _1158_ = sel_i[2] ? _1157_ : _1156_;
  assign _1159_ = sel_i[1] ? _0427_ : _0428_;
  assign _1160_ = sel_i[1] ? _0430_ : _0431_;
  assign _1161_ = sel_i[2] ? _1160_ : _1159_;
  assign _1162_ = sel_i[3] ? _1161_ : _1158_;
  assign _1163_ = sel_i[1] ? _0435_ : _0436_;
  assign _1164_ = sel_i[1] ? _0438_ : _0439_;
  assign _1165_ = sel_i[2] ? _1164_ : _1163_;
  assign _1166_ = sel_i[1] ? _0442_ : _0443_;
  assign _1167_ = sel_i[1] ? _0445_ : _0446_;
  assign _1168_ = sel_i[2] ? _1167_ : _1166_;
  assign _1169_ = sel_i[3] ? _1168_ : _1165_;
  assign data_o[46] = sel_i[4] ? _1169_ : _1162_;
  assign _1170_ = sel_i[1] ? _0450_ : _0451_;
  assign _1171_ = sel_i[1] ? _0453_ : _0454_;
  assign _1172_ = sel_i[2] ? _1171_ : _1170_;
  assign _1173_ = sel_i[1] ? _0457_ : _0458_;
  assign _1174_ = sel_i[1] ? _0460_ : _0461_;
  assign _1175_ = sel_i[2] ? _1174_ : _1173_;
  assign _1176_ = sel_i[3] ? _1175_ : _1172_;
  assign _1177_ = sel_i[1] ? _0465_ : _0466_;
  assign _1178_ = sel_i[1] ? _0468_ : _0469_;
  assign _1179_ = sel_i[2] ? _1178_ : _1177_;
  assign _1180_ = sel_i[1] ? _0472_ : _0473_;
  assign _1181_ = sel_i[1] ? _0475_ : _0476_;
  assign _1182_ = sel_i[2] ? _1181_ : _1180_;
  assign _1183_ = sel_i[3] ? _1182_ : _1179_;
  assign data_o[47] = sel_i[4] ? _1183_ : _1176_;
  assign _1184_ = sel_i[1] ? _0480_ : _0481_;
  assign _1185_ = sel_i[1] ? _0483_ : _0484_;
  assign _1186_ = sel_i[2] ? _1185_ : _1184_;
  assign _1187_ = sel_i[1] ? _0487_ : _0488_;
  assign _1188_ = sel_i[1] ? _0490_ : _0491_;
  assign _1189_ = sel_i[2] ? _1188_ : _1187_;
  assign _1190_ = sel_i[3] ? _1189_ : _1186_;
  assign _1191_ = sel_i[1] ? _0495_ : _0496_;
  assign _1192_ = sel_i[1] ? _0498_ : _0499_;
  assign _1193_ = sel_i[2] ? _1192_ : _1191_;
  assign _1194_ = sel_i[1] ? _0502_ : _0503_;
  assign _1195_ = sel_i[1] ? _0505_ : _0506_;
  assign _1196_ = sel_i[2] ? _1195_ : _1194_;
  assign _1197_ = sel_i[3] ? _1196_ : _1193_;
  assign data_o[48] = sel_i[4] ? _1197_ : _1190_;
  assign _1198_ = sel_i[1] ? _0510_ : _0511_;
  assign _1199_ = sel_i[1] ? _0513_ : _0514_;
  assign _1200_ = sel_i[2] ? _1199_ : _1198_;
  assign _1201_ = sel_i[1] ? _0517_ : _0518_;
  assign _1202_ = sel_i[1] ? _0520_ : _0521_;
  assign _1203_ = sel_i[2] ? _1202_ : _1201_;
  assign _1204_ = sel_i[3] ? _1203_ : _1200_;
  assign _1205_ = sel_i[1] ? _0525_ : _0526_;
  assign _1206_ = sel_i[1] ? _0528_ : _0529_;
  assign _1207_ = sel_i[2] ? _1206_ : _1205_;
  assign _1208_ = sel_i[1] ? _0532_ : _0533_;
  assign _1209_ = sel_i[1] ? _0535_ : _0536_;
  assign _1210_ = sel_i[2] ? _1209_ : _1208_;
  assign _1211_ = sel_i[3] ? _1210_ : _1207_;
  assign data_o[49] = sel_i[4] ? _1211_ : _1204_;
  assign _1212_ = sel_i[1] ? _0540_ : _0541_;
  assign _1213_ = sel_i[1] ? _0543_ : _0544_;
  assign _1214_ = sel_i[2] ? _1213_ : _1212_;
  assign _1215_ = sel_i[1] ? _0547_ : _0548_;
  assign _1216_ = sel_i[1] ? _0550_ : _0551_;
  assign _1217_ = sel_i[2] ? _1216_ : _1215_;
  assign _1218_ = sel_i[3] ? _1217_ : _1214_;
  assign _1219_ = sel_i[1] ? _0555_ : _0556_;
  assign _1220_ = sel_i[1] ? _0558_ : _0559_;
  assign _1221_ = sel_i[2] ? _1220_ : _1219_;
  assign _1222_ = sel_i[1] ? _0562_ : _0563_;
  assign _1223_ = sel_i[1] ? _0565_ : _0566_;
  assign _1224_ = sel_i[2] ? _1223_ : _1222_;
  assign _1225_ = sel_i[3] ? _1224_ : _1221_;
  assign data_o[50] = sel_i[4] ? _1225_ : _1218_;
  assign _1226_ = sel_i[1] ? _0570_ : _0571_;
  assign _1227_ = sel_i[1] ? _0573_ : _0574_;
  assign _1228_ = sel_i[2] ? _1227_ : _1226_;
  assign _1229_ = sel_i[1] ? _0577_ : _0578_;
  assign _1230_ = sel_i[1] ? _0580_ : _0581_;
  assign _1231_ = sel_i[2] ? _1230_ : _1229_;
  assign _1232_ = sel_i[3] ? _1231_ : _1228_;
  assign _1233_ = sel_i[1] ? _0585_ : _0586_;
  assign _1234_ = sel_i[1] ? _0588_ : _0589_;
  assign _1235_ = sel_i[2] ? _1234_ : _1233_;
  assign _1236_ = sel_i[1] ? _0592_ : _0593_;
  assign _1237_ = sel_i[1] ? _0595_ : _0596_;
  assign _1238_ = sel_i[2] ? _1237_ : _1236_;
  assign _1239_ = sel_i[3] ? _1238_ : _1235_;
  assign data_o[51] = sel_i[4] ? _1239_ : _1232_;
  assign _1240_ = sel_i[1] ? _0600_ : _0601_;
  assign _1241_ = sel_i[1] ? _0603_ : _0604_;
  assign _1242_ = sel_i[2] ? _1241_ : _1240_;
  assign _1243_ = sel_i[1] ? _0607_ : _0608_;
  assign _1244_ = sel_i[1] ? _0610_ : _0611_;
  assign _1245_ = sel_i[2] ? _1244_ : _1243_;
  assign _1246_ = sel_i[3] ? _1245_ : _1242_;
  assign _1247_ = sel_i[1] ? _0615_ : _0616_;
  assign _1248_ = sel_i[1] ? _0618_ : _0619_;
  assign _1249_ = sel_i[2] ? _1248_ : _1247_;
  assign _1250_ = sel_i[1] ? _0622_ : _0623_;
  assign _1251_ = sel_i[1] ? _0625_ : _0626_;
  assign _1252_ = sel_i[2] ? _1251_ : _1250_;
  assign _1253_ = sel_i[3] ? _1252_ : _1249_;
  assign data_o[52] = sel_i[4] ? _1253_ : _1246_;
  assign _1254_ = sel_i[1] ? _0630_ : _0631_;
  assign _1255_ = sel_i[1] ? _0633_ : _0634_;
  assign _1256_ = sel_i[2] ? _1255_ : _1254_;
  assign _1257_ = sel_i[1] ? _0637_ : _0638_;
  assign _1258_ = sel_i[1] ? _0640_ : _0641_;
  assign _1259_ = sel_i[2] ? _1258_ : _1257_;
  assign _1260_ = sel_i[3] ? _1259_ : _1256_;
  assign _1261_ = sel_i[1] ? _0645_ : _0646_;
  assign _1262_ = sel_i[1] ? _0648_ : _0649_;
  assign _1263_ = sel_i[2] ? _1262_ : _1261_;
  assign _1264_ = sel_i[1] ? _0652_ : _0653_;
  assign _1265_ = sel_i[1] ? _0655_ : _0656_;
  assign _1266_ = sel_i[2] ? _1265_ : _1264_;
  assign _1267_ = sel_i[3] ? _1266_ : _1263_;
  assign data_o[53] = sel_i[4] ? _1267_ : _1260_;
  assign _1268_ = sel_i[1] ? _0660_ : _0661_;
  assign _1269_ = sel_i[1] ? _0663_ : _0664_;
  assign _1270_ = sel_i[2] ? _1269_ : _1268_;
  assign _1271_ = sel_i[1] ? _0667_ : _0668_;
  assign _1272_ = sel_i[1] ? _0670_ : _0671_;
  assign _1273_ = sel_i[2] ? _1272_ : _1271_;
  assign _1274_ = sel_i[3] ? _1273_ : _1270_;
  assign _1275_ = sel_i[1] ? _0675_ : _0676_;
  assign _1276_ = sel_i[1] ? _0678_ : _0679_;
  assign _1277_ = sel_i[2] ? _1276_ : _1275_;
  assign _1278_ = sel_i[1] ? _0682_ : _0683_;
  assign _1279_ = sel_i[1] ? _0685_ : _0686_;
  assign _1280_ = sel_i[2] ? _1279_ : _1278_;
  assign _1281_ = sel_i[3] ? _1280_ : _1277_;
  assign data_o[54] = sel_i[4] ? _1281_ : _1274_;
  assign _1282_ = sel_i[1] ? _0690_ : _0691_;
  assign _1283_ = sel_i[1] ? _0693_ : _0694_;
  assign _1284_ = sel_i[2] ? _1283_ : _1282_;
  assign _1285_ = sel_i[1] ? _0697_ : _0698_;
  assign _1286_ = sel_i[1] ? _0700_ : _0701_;
  assign _1287_ = sel_i[2] ? _1286_ : _1285_;
  assign _1288_ = sel_i[3] ? _1287_ : _1284_;
  assign _1289_ = sel_i[1] ? _0705_ : _0706_;
  assign _1290_ = sel_i[1] ? _0708_ : _0709_;
  assign _1291_ = sel_i[2] ? _1290_ : _1289_;
  assign _1292_ = sel_i[1] ? _0712_ : _0713_;
  assign _1293_ = sel_i[1] ? _0715_ : _0716_;
  assign _1294_ = sel_i[2] ? _1293_ : _1292_;
  assign _1295_ = sel_i[3] ? _1294_ : _1291_;
  assign data_o[55] = sel_i[4] ? _1295_ : _1288_;
  assign _1296_ = sel_i[1] ? _0720_ : _0721_;
  assign _1297_ = sel_i[1] ? _0723_ : _0724_;
  assign _1298_ = sel_i[2] ? _1297_ : _1296_;
  assign _1299_ = sel_i[1] ? _0727_ : _0728_;
  assign _1300_ = sel_i[1] ? _0730_ : _0731_;
  assign _1301_ = sel_i[2] ? _1300_ : _1299_;
  assign _1302_ = sel_i[3] ? _1301_ : _1298_;
  assign _1303_ = sel_i[1] ? _0735_ : _0736_;
  assign _1304_ = sel_i[1] ? _0738_ : _0739_;
  assign _1305_ = sel_i[2] ? _1304_ : _1303_;
  assign _1306_ = sel_i[1] ? _0742_ : _0743_;
  assign _1307_ = sel_i[1] ? _0745_ : _0746_;
  assign _1308_ = sel_i[2] ? _1307_ : _1306_;
  assign _1309_ = sel_i[3] ? _1308_ : _1305_;
  assign data_o[56] = sel_i[4] ? _1309_ : _1302_;
  assign _1310_ = sel_i[1] ? _0750_ : _0751_;
  assign _1311_ = sel_i[1] ? _0753_ : _0754_;
  assign _1312_ = sel_i[2] ? _1311_ : _1310_;
  assign _1313_ = sel_i[1] ? _0757_ : _0758_;
  assign _1314_ = sel_i[1] ? _0760_ : _0761_;
  assign _1315_ = sel_i[2] ? _1314_ : _1313_;
  assign _1316_ = sel_i[3] ? _1315_ : _1312_;
  assign _1317_ = sel_i[1] ? _0765_ : _0766_;
  assign _1318_ = sel_i[1] ? _0768_ : _0769_;
  assign _1319_ = sel_i[2] ? _1318_ : _1317_;
  assign _1320_ = sel_i[1] ? _0772_ : _0773_;
  assign _1321_ = sel_i[1] ? _0775_ : _0776_;
  assign _1322_ = sel_i[2] ? _1321_ : _1320_;
  assign _1323_ = sel_i[3] ? _1322_ : _1319_;
  assign data_o[57] = sel_i[4] ? _1323_ : _1316_;
  assign _1324_ = sel_i[1] ? _0780_ : _0781_;
  assign _1325_ = sel_i[1] ? _0783_ : _0784_;
  assign _1326_ = sel_i[2] ? _1325_ : _1324_;
  assign _1327_ = sel_i[1] ? _0787_ : _0788_;
  assign _1328_ = sel_i[1] ? _0790_ : _0791_;
  assign _1329_ = sel_i[2] ? _1328_ : _1327_;
  assign _1330_ = sel_i[3] ? _1329_ : _1326_;
  assign _1331_ = sel_i[1] ? _0795_ : _0796_;
  assign _1332_ = sel_i[1] ? _0798_ : _0799_;
  assign _1333_ = sel_i[2] ? _1332_ : _1331_;
  assign _1334_ = sel_i[1] ? _0802_ : _0803_;
  assign _1335_ = sel_i[1] ? _0805_ : _0806_;
  assign _1336_ = sel_i[2] ? _1335_ : _1334_;
  assign _1337_ = sel_i[3] ? _1336_ : _1333_;
  assign data_o[58] = sel_i[4] ? _1337_ : _1330_;
  assign _1338_ = sel_i[1] ? _0810_ : _0811_;
  assign _1339_ = sel_i[1] ? _0813_ : _0814_;
  assign _1340_ = sel_i[2] ? _1339_ : _1338_;
  assign _1341_ = sel_i[1] ? _0817_ : _0818_;
  assign _1342_ = sel_i[1] ? _0820_ : _0821_;
  assign _1343_ = sel_i[2] ? _1342_ : _1341_;
  assign _1344_ = sel_i[3] ? _1343_ : _1340_;
  assign _1345_ = sel_i[1] ? _0825_ : _0826_;
  assign _1346_ = sel_i[1] ? _0828_ : _0829_;
  assign _1347_ = sel_i[2] ? _1346_ : _1345_;
  assign _1348_ = sel_i[1] ? _0832_ : _0833_;
  assign _1349_ = sel_i[1] ? _0835_ : _0836_;
  assign _1350_ = sel_i[2] ? _1349_ : _1348_;
  assign _1351_ = sel_i[3] ? _1350_ : _1347_;
  assign data_o[59] = sel_i[4] ? _1351_ : _1344_;
  assign _1352_ = sel_i[1] ? _0840_ : _0841_;
  assign _1353_ = sel_i[1] ? _0843_ : _0844_;
  assign _1354_ = sel_i[2] ? _1353_ : _1352_;
  assign _1355_ = sel_i[1] ? _0847_ : _0848_;
  assign _1356_ = sel_i[1] ? _0850_ : _0851_;
  assign _1357_ = sel_i[2] ? _1356_ : _1355_;
  assign _1358_ = sel_i[3] ? _1357_ : _1354_;
  assign _1359_ = sel_i[1] ? _0855_ : _0856_;
  assign _1360_ = sel_i[1] ? _0858_ : _0859_;
  assign _1361_ = sel_i[2] ? _1360_ : _1359_;
  assign _1362_ = sel_i[1] ? _0862_ : _0863_;
  assign _1363_ = sel_i[1] ? _0865_ : _0866_;
  assign _1364_ = sel_i[2] ? _1363_ : _1362_;
  assign _1365_ = sel_i[3] ? _1364_ : _1361_;
  assign data_o[60] = sel_i[4] ? _1365_ : _1358_;
  assign _1366_ = sel_i[1] ? _0870_ : _0871_;
  assign _1367_ = sel_i[1] ? _0873_ : _0874_;
  assign _1368_ = sel_i[2] ? _1367_ : _1366_;
  assign _1369_ = sel_i[1] ? _0877_ : _0878_;
  assign _1370_ = sel_i[1] ? _0880_ : _0881_;
  assign _1371_ = sel_i[2] ? _1370_ : _1369_;
  assign _1372_ = sel_i[3] ? _1371_ : _1368_;
  assign _1373_ = sel_i[1] ? _0885_ : _0886_;
  assign _1374_ = sel_i[1] ? _0888_ : _0889_;
  assign _1375_ = sel_i[2] ? _1374_ : _1373_;
  assign _1376_ = sel_i[1] ? _0892_ : _0893_;
  assign _1377_ = sel_i[1] ? _0895_ : _0896_;
  assign _1378_ = sel_i[2] ? _1377_ : _1376_;
  assign _1379_ = sel_i[3] ? _1378_ : _1375_;
  assign data_o[61] = sel_i[4] ? _1379_ : _1372_;
  assign _1380_ = sel_i[1] ? _0900_ : _0901_;
  assign _1381_ = sel_i[1] ? _0903_ : _0904_;
  assign _1382_ = sel_i[2] ? _1381_ : _1380_;
  assign _1383_ = sel_i[1] ? _0907_ : _0908_;
  assign _1384_ = sel_i[1] ? _0910_ : _0911_;
  assign _1385_ = sel_i[2] ? _1384_ : _1383_;
  assign _1386_ = sel_i[3] ? _1385_ : _1382_;
  assign _1387_ = sel_i[1] ? _0915_ : _0916_;
  assign _1388_ = sel_i[1] ? _0918_ : _0919_;
  assign _1389_ = sel_i[2] ? _1388_ : _1387_;
  assign _1390_ = sel_i[1] ? _0922_ : _0923_;
  assign _1391_ = sel_i[1] ? _0925_ : _0926_;
  assign _1392_ = sel_i[2] ? _1391_ : _1390_;
  assign _1393_ = sel_i[3] ? _1392_ : _1389_;
  assign data_o[62] = sel_i[4] ? _1393_ : _1386_;
  assign _1394_ = sel_i[1] ? _0930_ : _0931_;
  assign _1395_ = sel_i[1] ? _0933_ : _0934_;
  assign _1396_ = sel_i[2] ? _1395_ : _1394_;
  assign _1397_ = sel_i[1] ? _0937_ : _0938_;
  assign _1398_ = sel_i[1] ? _0940_ : _0941_;
  assign _1399_ = sel_i[2] ? _1398_ : _1397_;
  assign _1400_ = sel_i[3] ? _1399_ : _1396_;
  assign _1401_ = sel_i[1] ? _0945_ : _0946_;
  assign _1402_ = sel_i[1] ? _0948_ : _0949_;
  assign _1403_ = sel_i[2] ? _1402_ : _1401_;
  assign _1404_ = sel_i[1] ? _0952_ : _0953_;
  assign _1405_ = sel_i[1] ? _0955_ : _0956_;
  assign _1406_ = sel_i[2] ? _1405_ : _1404_;
  assign _1407_ = sel_i[3] ? _1406_ : _1403_;
  assign data_o[63] = sel_i[4] ? _1407_ : _1400_;
  assign _1408_ = sel_i[2] ? _0002_ : _0005_;
  assign _1409_ = sel_i[2] ? _0009_ : _0012_;
  assign _1410_ = sel_i[3] ? _1409_ : _1408_;
  assign _1411_ = sel_i[2] ? _0017_ : _0020_;
  assign _1412_ = sel_i[2] ? _0024_ : _0027_;
  assign _1413_ = sel_i[3] ? _1412_ : _1411_;
  assign data_o[64] = sel_i[4] ? _1413_ : _1410_;
  assign _1414_ = sel_i[2] ? _0032_ : _0035_;
  assign _1415_ = sel_i[2] ? _0039_ : _0042_;
  assign _1416_ = sel_i[3] ? _1415_ : _1414_;
  assign _1417_ = sel_i[2] ? _0047_ : _0050_;
  assign _1418_ = sel_i[2] ? _0054_ : _0057_;
  assign _1419_ = sel_i[3] ? _1418_ : _1417_;
  assign data_o[65] = sel_i[4] ? _1419_ : _1416_;
  assign _1420_ = sel_i[2] ? _0062_ : _0065_;
  assign _1421_ = sel_i[2] ? _0069_ : _0072_;
  assign _1422_ = sel_i[3] ? _1421_ : _1420_;
  assign _1423_ = sel_i[2] ? _0077_ : _0080_;
  assign _1424_ = sel_i[2] ? _0084_ : _0087_;
  assign _1425_ = sel_i[3] ? _1424_ : _1423_;
  assign data_o[66] = sel_i[4] ? _1425_ : _1422_;
  assign _1426_ = sel_i[2] ? _0092_ : _0095_;
  assign _1427_ = sel_i[2] ? _0099_ : _0102_;
  assign _1428_ = sel_i[3] ? _1427_ : _1426_;
  assign _1429_ = sel_i[2] ? _0107_ : _0110_;
  assign _1430_ = sel_i[2] ? _0114_ : _0117_;
  assign _1431_ = sel_i[3] ? _1430_ : _1429_;
  assign data_o[67] = sel_i[4] ? _1431_ : _1428_;
  assign _1432_ = sel_i[2] ? _0122_ : _0125_;
  assign _1433_ = sel_i[2] ? _0129_ : _0132_;
  assign _1434_ = sel_i[3] ? _1433_ : _1432_;
  assign _1435_ = sel_i[2] ? _0137_ : _0140_;
  assign _1436_ = sel_i[2] ? _0144_ : _0147_;
  assign _1437_ = sel_i[3] ? _1436_ : _1435_;
  assign data_o[68] = sel_i[4] ? _1437_ : _1434_;
  assign _1438_ = sel_i[2] ? _0152_ : _0155_;
  assign _1439_ = sel_i[2] ? _0159_ : _0162_;
  assign _1440_ = sel_i[3] ? _1439_ : _1438_;
  assign _1441_ = sel_i[2] ? _0167_ : _0170_;
  assign _1442_ = sel_i[2] ? _0174_ : _0177_;
  assign _1443_ = sel_i[3] ? _1442_ : _1441_;
  assign data_o[69] = sel_i[4] ? _1443_ : _1440_;
  assign _1444_ = sel_i[2] ? _0182_ : _0185_;
  assign _1445_ = sel_i[2] ? _0189_ : _0192_;
  assign _1446_ = sel_i[3] ? _1445_ : _1444_;
  assign _1447_ = sel_i[2] ? _0197_ : _0200_;
  assign _1448_ = sel_i[2] ? _0204_ : _0207_;
  assign _1449_ = sel_i[3] ? _1448_ : _1447_;
  assign data_o[70] = sel_i[4] ? _1449_ : _1446_;
  assign _1450_ = sel_i[2] ? _0212_ : _0215_;
  assign _1451_ = sel_i[2] ? _0219_ : _0222_;
  assign _1452_ = sel_i[3] ? _1451_ : _1450_;
  assign _1453_ = sel_i[2] ? _0227_ : _0230_;
  assign _1454_ = sel_i[2] ? _0234_ : _0237_;
  assign _1455_ = sel_i[3] ? _1454_ : _1453_;
  assign data_o[71] = sel_i[4] ? _1455_ : _1452_;
  assign _1456_ = sel_i[2] ? _0242_ : _0245_;
  assign _1457_ = sel_i[2] ? _0249_ : _0252_;
  assign _1458_ = sel_i[3] ? _1457_ : _1456_;
  assign _1459_ = sel_i[2] ? _0257_ : _0260_;
  assign _1460_ = sel_i[2] ? _0264_ : _0267_;
  assign _1461_ = sel_i[3] ? _1460_ : _1459_;
  assign data_o[72] = sel_i[4] ? _1461_ : _1458_;
  assign _1462_ = sel_i[2] ? _0272_ : _0275_;
  assign _1463_ = sel_i[2] ? _0279_ : _0282_;
  assign _1464_ = sel_i[3] ? _1463_ : _1462_;
  assign _1465_ = sel_i[2] ? _0287_ : _0290_;
  assign _1466_ = sel_i[2] ? _0294_ : _0297_;
  assign _1467_ = sel_i[3] ? _1466_ : _1465_;
  assign data_o[73] = sel_i[4] ? _1467_ : _1464_;
  assign _1468_ = sel_i[2] ? _0302_ : _0305_;
  assign _1469_ = sel_i[2] ? _0309_ : _0312_;
  assign _1470_ = sel_i[3] ? _1469_ : _1468_;
  assign _1471_ = sel_i[2] ? _0317_ : _0320_;
  assign _1472_ = sel_i[2] ? _0324_ : _0327_;
  assign _1473_ = sel_i[3] ? _1472_ : _1471_;
  assign data_o[74] = sel_i[4] ? _1473_ : _1470_;
  assign _1474_ = sel_i[2] ? _0332_ : _0335_;
  assign _1475_ = sel_i[2] ? _0339_ : _0342_;
  assign _1476_ = sel_i[3] ? _1475_ : _1474_;
  assign _1477_ = sel_i[2] ? _0347_ : _0350_;
  assign _1478_ = sel_i[2] ? _0354_ : _0357_;
  assign _1479_ = sel_i[3] ? _1478_ : _1477_;
  assign data_o[75] = sel_i[4] ? _1479_ : _1476_;
  assign _1480_ = sel_i[2] ? _0362_ : _0365_;
  assign _1481_ = sel_i[2] ? _0369_ : _0372_;
  assign _1482_ = sel_i[3] ? _1481_ : _1480_;
  assign _1483_ = sel_i[2] ? _0377_ : _0380_;
  assign _1484_ = sel_i[2] ? _0384_ : _0387_;
  assign _1485_ = sel_i[3] ? _1484_ : _1483_;
  assign data_o[76] = sel_i[4] ? _1485_ : _1482_;
  assign _1486_ = sel_i[2] ? _0392_ : _0395_;
  assign _1487_ = sel_i[2] ? _0399_ : _0402_;
  assign _1488_ = sel_i[3] ? _1487_ : _1486_;
  assign _1489_ = sel_i[2] ? _0407_ : _0410_;
  assign _1490_ = sel_i[2] ? _0414_ : _0417_;
  assign _1491_ = sel_i[3] ? _1490_ : _1489_;
  assign data_o[77] = sel_i[4] ? _1491_ : _1488_;
  assign _1492_ = sel_i[2] ? _0422_ : _0425_;
  assign _1493_ = sel_i[2] ? _0429_ : _0432_;
  assign _1494_ = sel_i[3] ? _1493_ : _1492_;
  assign _1495_ = sel_i[2] ? _0437_ : _0440_;
  assign _1496_ = sel_i[2] ? _0444_ : _0447_;
  assign _1497_ = sel_i[3] ? _1496_ : _1495_;
  assign data_o[78] = sel_i[4] ? _1497_ : _1494_;
  assign _1498_ = sel_i[2] ? _0452_ : _0455_;
  assign _1499_ = sel_i[2] ? _0459_ : _0462_;
  assign _1500_ = sel_i[3] ? _1499_ : _1498_;
  assign _1501_ = sel_i[2] ? _0467_ : _0470_;
  assign _1502_ = sel_i[2] ? _0474_ : _0477_;
  assign _1503_ = sel_i[3] ? _1502_ : _1501_;
  assign data_o[79] = sel_i[4] ? _1503_ : _1500_;
  assign _1504_ = sel_i[2] ? _0482_ : _0485_;
  assign _1505_ = sel_i[2] ? _0489_ : _0492_;
  assign _1506_ = sel_i[3] ? _1505_ : _1504_;
  assign _1507_ = sel_i[2] ? _0497_ : _0500_;
  assign _1508_ = sel_i[2] ? _0504_ : _0507_;
  assign _1509_ = sel_i[3] ? _1508_ : _1507_;
  assign data_o[80] = sel_i[4] ? _1509_ : _1506_;
  assign _1510_ = sel_i[2] ? _0512_ : _0515_;
  assign _1511_ = sel_i[2] ? _0519_ : _0522_;
  assign _1512_ = sel_i[3] ? _1511_ : _1510_;
  assign _1513_ = sel_i[2] ? _0527_ : _0530_;
  assign _1514_ = sel_i[2] ? _0534_ : _0537_;
  assign _1515_ = sel_i[3] ? _1514_ : _1513_;
  assign data_o[81] = sel_i[4] ? _1515_ : _1512_;
  assign _1516_ = sel_i[2] ? _0542_ : _0545_;
  assign _1517_ = sel_i[2] ? _0549_ : _0552_;
  assign _1518_ = sel_i[3] ? _1517_ : _1516_;
  assign _1519_ = sel_i[2] ? _0557_ : _0560_;
  assign _1520_ = sel_i[2] ? _0564_ : _0567_;
  assign _1521_ = sel_i[3] ? _1520_ : _1519_;
  assign data_o[82] = sel_i[4] ? _1521_ : _1518_;
  assign _1522_ = sel_i[2] ? _0572_ : _0575_;
  assign _1523_ = sel_i[2] ? _0579_ : _0582_;
  assign _1524_ = sel_i[3] ? _1523_ : _1522_;
  assign _1525_ = sel_i[2] ? _0587_ : _0590_;
  assign _1526_ = sel_i[2] ? _0594_ : _0597_;
  assign _1527_ = sel_i[3] ? _1526_ : _1525_;
  assign data_o[83] = sel_i[4] ? _1527_ : _1524_;
  assign _1528_ = sel_i[2] ? _0602_ : _0605_;
  assign _1529_ = sel_i[2] ? _0609_ : _0612_;
  assign _1530_ = sel_i[3] ? _1529_ : _1528_;
  assign _1531_ = sel_i[2] ? _0617_ : _0620_;
  assign _1532_ = sel_i[2] ? _0624_ : _0627_;
  assign _1533_ = sel_i[3] ? _1532_ : _1531_;
  assign data_o[84] = sel_i[4] ? _1533_ : _1530_;
  assign _1534_ = sel_i[2] ? _0632_ : _0635_;
  assign _1535_ = sel_i[2] ? _0639_ : _0642_;
  assign _1536_ = sel_i[3] ? _1535_ : _1534_;
  assign _1537_ = sel_i[2] ? _0647_ : _0650_;
  assign _1538_ = sel_i[2] ? _0654_ : _0657_;
  assign _1539_ = sel_i[3] ? _1538_ : _1537_;
  assign data_o[85] = sel_i[4] ? _1539_ : _1536_;
  assign _1540_ = sel_i[2] ? _0662_ : _0665_;
  assign _1541_ = sel_i[2] ? _0669_ : _0672_;
  assign _1542_ = sel_i[3] ? _1541_ : _1540_;
  assign _1543_ = sel_i[2] ? _0677_ : _0680_;
  assign _1544_ = sel_i[2] ? _0684_ : _0687_;
  assign _1545_ = sel_i[3] ? _1544_ : _1543_;
  assign data_o[86] = sel_i[4] ? _1545_ : _1542_;
  assign _1546_ = sel_i[2] ? _0692_ : _0695_;
  assign _1547_ = sel_i[2] ? _0699_ : _0702_;
  assign _1548_ = sel_i[3] ? _1547_ : _1546_;
  assign _1549_ = sel_i[2] ? _0707_ : _0710_;
  assign _1550_ = sel_i[2] ? _0714_ : _0717_;
  assign _1551_ = sel_i[3] ? _1550_ : _1549_;
  assign data_o[87] = sel_i[4] ? _1551_ : _1548_;
  assign _1552_ = sel_i[2] ? _0722_ : _0725_;
  assign _1553_ = sel_i[2] ? _0729_ : _0732_;
  assign _1554_ = sel_i[3] ? _1553_ : _1552_;
  assign _1555_ = sel_i[2] ? _0737_ : _0740_;
  assign _1556_ = sel_i[2] ? _0744_ : _0747_;
  assign _1557_ = sel_i[3] ? _1556_ : _1555_;
  assign data_o[88] = sel_i[4] ? _1557_ : _1554_;
  assign _1558_ = sel_i[2] ? _0752_ : _0755_;
  assign _1559_ = sel_i[2] ? _0759_ : _0762_;
  assign _1560_ = sel_i[3] ? _1559_ : _1558_;
  assign _1561_ = sel_i[2] ? _0767_ : _0770_;
  assign _1562_ = sel_i[2] ? _0774_ : _0777_;
  assign _1563_ = sel_i[3] ? _1562_ : _1561_;
  assign data_o[89] = sel_i[4] ? _1563_ : _1560_;
  assign _1564_ = sel_i[2] ? _0782_ : _0785_;
  assign _1565_ = sel_i[2] ? _0789_ : _0792_;
  assign _1566_ = sel_i[3] ? _1565_ : _1564_;
  assign _1567_ = sel_i[2] ? _0797_ : _0800_;
  assign _1568_ = sel_i[2] ? _0804_ : _0807_;
  assign _1569_ = sel_i[3] ? _1568_ : _1567_;
  assign data_o[90] = sel_i[4] ? _1569_ : _1566_;
  assign _1570_ = sel_i[2] ? _0812_ : _0815_;
  assign _1571_ = sel_i[2] ? _0819_ : _0822_;
  assign _1572_ = sel_i[3] ? _1571_ : _1570_;
  assign _1573_ = sel_i[2] ? _0827_ : _0830_;
  assign _1574_ = sel_i[2] ? _0834_ : _0837_;
  assign _1575_ = sel_i[3] ? _1574_ : _1573_;
  assign data_o[91] = sel_i[4] ? _1575_ : _1572_;
  assign _1576_ = sel_i[2] ? _0842_ : _0845_;
  assign _1577_ = sel_i[2] ? _0849_ : _0852_;
  assign _1578_ = sel_i[3] ? _1577_ : _1576_;
  assign _1579_ = sel_i[2] ? _0857_ : _0860_;
  assign _1580_ = sel_i[2] ? _0864_ : _0867_;
  assign _1581_ = sel_i[3] ? _1580_ : _1579_;
  assign data_o[92] = sel_i[4] ? _1581_ : _1578_;
  assign _1582_ = sel_i[2] ? _0872_ : _0875_;
  assign _1583_ = sel_i[2] ? _0879_ : _0882_;
  assign _1584_ = sel_i[3] ? _1583_ : _1582_;
  assign _1585_ = sel_i[2] ? _0887_ : _0890_;
  assign _1586_ = sel_i[2] ? _0894_ : _0897_;
  assign _1587_ = sel_i[3] ? _1586_ : _1585_;
  assign data_o[93] = sel_i[4] ? _1587_ : _1584_;
  assign _1588_ = sel_i[2] ? _0902_ : _0905_;
  assign _1589_ = sel_i[2] ? _0909_ : _0912_;
  assign _1590_ = sel_i[3] ? _1589_ : _1588_;
  assign _1591_ = sel_i[2] ? _0917_ : _0920_;
  assign _1592_ = sel_i[2] ? _0924_ : _0927_;
  assign _1593_ = sel_i[3] ? _1592_ : _1591_;
  assign data_o[94] = sel_i[4] ? _1593_ : _1590_;
  assign _1594_ = sel_i[2] ? _0932_ : _0935_;
  assign _1595_ = sel_i[2] ? _0939_ : _0942_;
  assign _1596_ = sel_i[3] ? _1595_ : _1594_;
  assign _1597_ = sel_i[2] ? _0947_ : _0950_;
  assign _1598_ = sel_i[2] ? _0954_ : _0957_;
  assign _1599_ = sel_i[3] ? _1598_ : _1597_;
  assign data_o[95] = sel_i[4] ? _1599_ : _1596_;
  assign _1600_ = sel_i[2] ? _0960_ : _0961_;
  assign _1601_ = sel_i[2] ? _0963_ : _0964_;
  assign _1602_ = sel_i[3] ? _1601_ : _1600_;
  assign _1603_ = sel_i[2] ? _0967_ : _0968_;
  assign _1604_ = sel_i[2] ? _0970_ : _0971_;
  assign _1605_ = sel_i[3] ? _1604_ : _1603_;
  assign data_o[96] = sel_i[4] ? _1605_ : _1602_;
  assign _1606_ = sel_i[2] ? _0974_ : _0975_;
  assign _1607_ = sel_i[2] ? _0977_ : _0978_;
  assign _1608_ = sel_i[3] ? _1607_ : _1606_;
  assign _1609_ = sel_i[2] ? _0981_ : _0982_;
  assign _1610_ = sel_i[2] ? _0984_ : _0985_;
  assign _1611_ = sel_i[3] ? _1610_ : _1609_;
  assign data_o[97] = sel_i[4] ? _1611_ : _1608_;
  assign _1612_ = sel_i[2] ? _0988_ : _0989_;
  assign _1613_ = sel_i[2] ? _0991_ : _0992_;
  assign _1614_ = sel_i[3] ? _1613_ : _1612_;
  assign _1615_ = sel_i[2] ? _0995_ : _0996_;
  assign _1616_ = sel_i[2] ? _0998_ : _0999_;
  assign _1617_ = sel_i[3] ? _1616_ : _1615_;
  assign data_o[98] = sel_i[4] ? _1617_ : _1614_;
  assign _1618_ = sel_i[2] ? _1002_ : _1003_;
  assign _1619_ = sel_i[2] ? _1005_ : _1006_;
  assign _1620_ = sel_i[3] ? _1619_ : _1618_;
  assign _1621_ = sel_i[2] ? _1009_ : _1010_;
  assign _1622_ = sel_i[2] ? _1012_ : _1013_;
  assign _1623_ = sel_i[3] ? _1622_ : _1621_;
  assign data_o[99] = sel_i[4] ? _1623_ : _1620_;
  assign _1624_ = sel_i[2] ? _1016_ : _1017_;
  assign _1625_ = sel_i[2] ? _1019_ : _1020_;
  assign _1626_ = sel_i[3] ? _1625_ : _1624_;
  assign _1627_ = sel_i[2] ? _1023_ : _1024_;
  assign _1628_ = sel_i[2] ? _1026_ : _1027_;
  assign _1629_ = sel_i[3] ? _1628_ : _1627_;
  assign data_o[100] = sel_i[4] ? _1629_ : _1626_;
  assign _1630_ = sel_i[2] ? _1030_ : _1031_;
  assign _1631_ = sel_i[2] ? _1033_ : _1034_;
  assign _1632_ = sel_i[3] ? _1631_ : _1630_;
  assign _1633_ = sel_i[2] ? _1037_ : _1038_;
  assign _1634_ = sel_i[2] ? _1040_ : _1041_;
  assign _1635_ = sel_i[3] ? _1634_ : _1633_;
  assign data_o[101] = sel_i[4] ? _1635_ : _1632_;
  assign _1636_ = sel_i[2] ? _1044_ : _1045_;
  assign _1637_ = sel_i[2] ? _1047_ : _1048_;
  assign _1638_ = sel_i[3] ? _1637_ : _1636_;
  assign _1639_ = sel_i[2] ? _1051_ : _1052_;
  assign _1640_ = sel_i[2] ? _1054_ : _1055_;
  assign _1641_ = sel_i[3] ? _1640_ : _1639_;
  assign data_o[102] = sel_i[4] ? _1641_ : _1638_;
  assign _1642_ = sel_i[2] ? _1058_ : _1059_;
  assign _1643_ = sel_i[2] ? _1061_ : _1062_;
  assign _1644_ = sel_i[3] ? _1643_ : _1642_;
  assign _1645_ = sel_i[2] ? _1065_ : _1066_;
  assign _1646_ = sel_i[2] ? _1068_ : _1069_;
  assign _1647_ = sel_i[3] ? _1646_ : _1645_;
  assign data_o[103] = sel_i[4] ? _1647_ : _1644_;
  assign _1648_ = sel_i[2] ? _1072_ : _1073_;
  assign _1649_ = sel_i[2] ? _1075_ : _1076_;
  assign _1650_ = sel_i[3] ? _1649_ : _1648_;
  assign _1651_ = sel_i[2] ? _1079_ : _1080_;
  assign _1652_ = sel_i[2] ? _1082_ : _1083_;
  assign _1653_ = sel_i[3] ? _1652_ : _1651_;
  assign data_o[104] = sel_i[4] ? _1653_ : _1650_;
  assign _1654_ = sel_i[2] ? _1086_ : _1087_;
  assign _1655_ = sel_i[2] ? _1089_ : _1090_;
  assign _1656_ = sel_i[3] ? _1655_ : _1654_;
  assign _1657_ = sel_i[2] ? _1093_ : _1094_;
  assign _1658_ = sel_i[2] ? _1096_ : _1097_;
  assign _1659_ = sel_i[3] ? _1658_ : _1657_;
  assign data_o[105] = sel_i[4] ? _1659_ : _1656_;
  assign _1660_ = sel_i[2] ? _1100_ : _1101_;
  assign _1661_ = sel_i[2] ? _1103_ : _1104_;
  assign _1662_ = sel_i[3] ? _1661_ : _1660_;
  assign _1663_ = sel_i[2] ? _1107_ : _1108_;
  assign _1664_ = sel_i[2] ? _1110_ : _1111_;
  assign _1665_ = sel_i[3] ? _1664_ : _1663_;
  assign data_o[106] = sel_i[4] ? _1665_ : _1662_;
  assign _1666_ = sel_i[2] ? _1114_ : _1115_;
  assign _1667_ = sel_i[2] ? _1117_ : _1118_;
  assign _1668_ = sel_i[3] ? _1667_ : _1666_;
  assign _1669_ = sel_i[2] ? _1121_ : _1122_;
  assign _1670_ = sel_i[2] ? _1124_ : _1125_;
  assign _1671_ = sel_i[3] ? _1670_ : _1669_;
  assign data_o[107] = sel_i[4] ? _1671_ : _1668_;
  assign _1672_ = sel_i[2] ? _1128_ : _1129_;
  assign _1673_ = sel_i[2] ? _1131_ : _1132_;
  assign _1674_ = sel_i[3] ? _1673_ : _1672_;
  assign _1675_ = sel_i[2] ? _1135_ : _1136_;
  assign _1676_ = sel_i[2] ? _1138_ : _1139_;
  assign _1677_ = sel_i[3] ? _1676_ : _1675_;
  assign data_o[108] = sel_i[4] ? _1677_ : _1674_;
  assign _1678_ = sel_i[2] ? _1142_ : _1143_;
  assign _1679_ = sel_i[2] ? _1145_ : _1146_;
  assign _1680_ = sel_i[3] ? _1679_ : _1678_;
  assign _1681_ = sel_i[2] ? _1149_ : _1150_;
  assign _1682_ = sel_i[2] ? _1152_ : _1153_;
  assign _1683_ = sel_i[3] ? _1682_ : _1681_;
  assign data_o[109] = sel_i[4] ? _1683_ : _1680_;
  assign _1684_ = sel_i[2] ? _1156_ : _1157_;
  assign _1685_ = sel_i[2] ? _1159_ : _1160_;
  assign _1686_ = sel_i[3] ? _1685_ : _1684_;
  assign _1687_ = sel_i[2] ? _1163_ : _1164_;
  assign _1688_ = sel_i[2] ? _1166_ : _1167_;
  assign _1689_ = sel_i[3] ? _1688_ : _1687_;
  assign data_o[110] = sel_i[4] ? _1689_ : _1686_;
  assign _1690_ = sel_i[2] ? _1170_ : _1171_;
  assign _1691_ = sel_i[2] ? _1173_ : _1174_;
  assign _1692_ = sel_i[3] ? _1691_ : _1690_;
  assign _1693_ = sel_i[2] ? _1177_ : _1178_;
  assign _1694_ = sel_i[2] ? _1180_ : _1181_;
  assign _1695_ = sel_i[3] ? _1694_ : _1693_;
  assign data_o[111] = sel_i[4] ? _1695_ : _1692_;
  assign _1696_ = sel_i[2] ? _1184_ : _1185_;
  assign _1697_ = sel_i[2] ? _1187_ : _1188_;
  assign _1698_ = sel_i[3] ? _1697_ : _1696_;
  assign _1699_ = sel_i[2] ? _1191_ : _1192_;
  assign _1700_ = sel_i[2] ? _1194_ : _1195_;
  assign _1701_ = sel_i[3] ? _1700_ : _1699_;
  assign data_o[112] = sel_i[4] ? _1701_ : _1698_;
  assign _1702_ = sel_i[2] ? _1198_ : _1199_;
  assign _1703_ = sel_i[2] ? _1201_ : _1202_;
  assign _1704_ = sel_i[3] ? _1703_ : _1702_;
  assign _1705_ = sel_i[2] ? _1205_ : _1206_;
  assign _1706_ = sel_i[2] ? _1208_ : _1209_;
  assign _1707_ = sel_i[3] ? _1706_ : _1705_;
  assign data_o[113] = sel_i[4] ? _1707_ : _1704_;
  assign _1708_ = sel_i[2] ? _1212_ : _1213_;
  assign _1709_ = sel_i[2] ? _1215_ : _1216_;
  assign _1710_ = sel_i[3] ? _1709_ : _1708_;
  assign _1711_ = sel_i[2] ? _1219_ : _1220_;
  assign _1712_ = sel_i[2] ? _1222_ : _1223_;
  assign _1713_ = sel_i[3] ? _1712_ : _1711_;
  assign data_o[114] = sel_i[4] ? _1713_ : _1710_;
  assign _1714_ = sel_i[2] ? _1226_ : _1227_;
  assign _1715_ = sel_i[2] ? _1229_ : _1230_;
  assign _1716_ = sel_i[3] ? _1715_ : _1714_;
  assign _1717_ = sel_i[2] ? _1233_ : _1234_;
  assign _1718_ = sel_i[2] ? _1236_ : _1237_;
  assign _1719_ = sel_i[3] ? _1718_ : _1717_;
  assign data_o[115] = sel_i[4] ? _1719_ : _1716_;
  assign _1720_ = sel_i[2] ? _1240_ : _1241_;
  assign _1721_ = sel_i[2] ? _1243_ : _1244_;
  assign _1722_ = sel_i[3] ? _1721_ : _1720_;
  assign _1723_ = sel_i[2] ? _1247_ : _1248_;
  assign _1724_ = sel_i[2] ? _1250_ : _1251_;
  assign _1725_ = sel_i[3] ? _1724_ : _1723_;
  assign data_o[116] = sel_i[4] ? _1725_ : _1722_;
  assign _1726_ = sel_i[2] ? _1254_ : _1255_;
  assign _1727_ = sel_i[2] ? _1257_ : _1258_;
  assign _1728_ = sel_i[3] ? _1727_ : _1726_;
  assign _1729_ = sel_i[2] ? _1261_ : _1262_;
  assign _1730_ = sel_i[2] ? _1264_ : _1265_;
  assign _1731_ = sel_i[3] ? _1730_ : _1729_;
  assign data_o[117] = sel_i[4] ? _1731_ : _1728_;
  assign _1732_ = sel_i[2] ? _1268_ : _1269_;
  assign _1733_ = sel_i[2] ? _1271_ : _1272_;
  assign _1734_ = sel_i[3] ? _1733_ : _1732_;
  assign _1735_ = sel_i[2] ? _1275_ : _1276_;
  assign _1736_ = sel_i[2] ? _1278_ : _1279_;
  assign _1737_ = sel_i[3] ? _1736_ : _1735_;
  assign data_o[118] = sel_i[4] ? _1737_ : _1734_;
  assign _1738_ = sel_i[2] ? _1282_ : _1283_;
  assign _1739_ = sel_i[2] ? _1285_ : _1286_;
  assign _1740_ = sel_i[3] ? _1739_ : _1738_;
  assign _1741_ = sel_i[2] ? _1289_ : _1290_;
  assign _1742_ = sel_i[2] ? _1292_ : _1293_;
  assign _1743_ = sel_i[3] ? _1742_ : _1741_;
  assign data_o[119] = sel_i[4] ? _1743_ : _1740_;
  assign _1744_ = sel_i[2] ? _1296_ : _1297_;
  assign _1745_ = sel_i[2] ? _1299_ : _1300_;
  assign _1746_ = sel_i[3] ? _1745_ : _1744_;
  assign _1747_ = sel_i[2] ? _1303_ : _1304_;
  assign _1748_ = sel_i[2] ? _1306_ : _1307_;
  assign _1749_ = sel_i[3] ? _1748_ : _1747_;
  assign data_o[120] = sel_i[4] ? _1749_ : _1746_;
  assign _1750_ = sel_i[2] ? _1310_ : _1311_;
  assign _1751_ = sel_i[2] ? _1313_ : _1314_;
  assign _1752_ = sel_i[3] ? _1751_ : _1750_;
  assign _1753_ = sel_i[2] ? _1317_ : _1318_;
  assign _1754_ = sel_i[2] ? _1320_ : _1321_;
  assign _1755_ = sel_i[3] ? _1754_ : _1753_;
  assign data_o[121] = sel_i[4] ? _1755_ : _1752_;
  assign _1756_ = sel_i[2] ? _1324_ : _1325_;
  assign _1757_ = sel_i[2] ? _1327_ : _1328_;
  assign _1758_ = sel_i[3] ? _1757_ : _1756_;
  assign _1759_ = sel_i[2] ? _1331_ : _1332_;
  assign _1760_ = sel_i[2] ? _1334_ : _1335_;
  assign _1761_ = sel_i[3] ? _1760_ : _1759_;
  assign data_o[122] = sel_i[4] ? _1761_ : _1758_;
  assign _1762_ = sel_i[2] ? _1338_ : _1339_;
  assign _1763_ = sel_i[2] ? _1341_ : _1342_;
  assign _1764_ = sel_i[3] ? _1763_ : _1762_;
  assign _1765_ = sel_i[2] ? _1345_ : _1346_;
  assign _1766_ = sel_i[2] ? _1348_ : _1349_;
  assign _1767_ = sel_i[3] ? _1766_ : _1765_;
  assign data_o[123] = sel_i[4] ? _1767_ : _1764_;
  assign _1768_ = sel_i[2] ? _1352_ : _1353_;
  assign _1769_ = sel_i[2] ? _1355_ : _1356_;
  assign _1770_ = sel_i[3] ? _1769_ : _1768_;
  assign _1771_ = sel_i[2] ? _1359_ : _1360_;
  assign _1772_ = sel_i[2] ? _1362_ : _1363_;
  assign _1773_ = sel_i[3] ? _1772_ : _1771_;
  assign data_o[124] = sel_i[4] ? _1773_ : _1770_;
  assign _1774_ = sel_i[2] ? _1366_ : _1367_;
  assign _1775_ = sel_i[2] ? _1369_ : _1370_;
  assign _1776_ = sel_i[3] ? _1775_ : _1774_;
  assign _1777_ = sel_i[2] ? _1373_ : _1374_;
  assign _1778_ = sel_i[2] ? _1376_ : _1377_;
  assign _1779_ = sel_i[3] ? _1778_ : _1777_;
  assign data_o[125] = sel_i[4] ? _1779_ : _1776_;
  assign _1780_ = sel_i[2] ? _1380_ : _1381_;
  assign _1781_ = sel_i[2] ? _1383_ : _1384_;
  assign _1782_ = sel_i[3] ? _1781_ : _1780_;
  assign _1783_ = sel_i[2] ? _1387_ : _1388_;
  assign _1784_ = sel_i[2] ? _1390_ : _1391_;
  assign _1785_ = sel_i[3] ? _1784_ : _1783_;
  assign data_o[126] = sel_i[4] ? _1785_ : _1782_;
  assign _1786_ = sel_i[2] ? _1394_ : _1395_;
  assign _1787_ = sel_i[2] ? _1397_ : _1398_;
  assign _1788_ = sel_i[3] ? _1787_ : _1786_;
  assign _1789_ = sel_i[2] ? _1401_ : _1402_;
  assign _1790_ = sel_i[2] ? _1404_ : _1405_;
  assign _1791_ = sel_i[3] ? _1790_ : _1789_;
  assign data_o[127] = sel_i[4] ? _1791_ : _1788_;
  assign _1792_ = sel_i[3] ? _0006_ : _0013_;
  assign _1793_ = sel_i[3] ? _0021_ : _0028_;
  assign data_o[128] = sel_i[4] ? _1793_ : _1792_;
  assign _1794_ = sel_i[3] ? _0036_ : _0043_;
  assign _1795_ = sel_i[3] ? _0051_ : _0058_;
  assign data_o[129] = sel_i[4] ? _1795_ : _1794_;
  assign _1796_ = sel_i[3] ? _0066_ : _0073_;
  assign _1797_ = sel_i[3] ? _0081_ : _0088_;
  assign data_o[130] = sel_i[4] ? _1797_ : _1796_;
  assign _1798_ = sel_i[3] ? _0096_ : _0103_;
  assign _1799_ = sel_i[3] ? _0111_ : _0118_;
  assign data_o[131] = sel_i[4] ? _1799_ : _1798_;
  assign _1800_ = sel_i[3] ? _0126_ : _0133_;
  assign _1801_ = sel_i[3] ? _0141_ : _0148_;
  assign data_o[132] = sel_i[4] ? _1801_ : _1800_;
  assign _1802_ = sel_i[3] ? _0156_ : _0163_;
  assign _1803_ = sel_i[3] ? _0171_ : _0178_;
  assign data_o[133] = sel_i[4] ? _1803_ : _1802_;
  assign _1804_ = sel_i[3] ? _0186_ : _0193_;
  assign _1805_ = sel_i[3] ? _0201_ : _0208_;
  assign data_o[134] = sel_i[4] ? _1805_ : _1804_;
  assign _1806_ = sel_i[3] ? _0216_ : _0223_;
  assign _1807_ = sel_i[3] ? _0231_ : _0238_;
  assign data_o[135] = sel_i[4] ? _1807_ : _1806_;
  assign _1808_ = sel_i[3] ? _0246_ : _0253_;
  assign _1809_ = sel_i[3] ? _0261_ : _0268_;
  assign data_o[136] = sel_i[4] ? _1809_ : _1808_;
  assign _1810_ = sel_i[3] ? _0276_ : _0283_;
  assign _1811_ = sel_i[3] ? _0291_ : _0298_;
  assign data_o[137] = sel_i[4] ? _1811_ : _1810_;
  assign _1812_ = sel_i[3] ? _0306_ : _0313_;
  assign _1813_ = sel_i[3] ? _0321_ : _0328_;
  assign data_o[138] = sel_i[4] ? _1813_ : _1812_;
  assign _1814_ = sel_i[3] ? _0336_ : _0343_;
  assign _1815_ = sel_i[3] ? _0351_ : _0358_;
  assign data_o[139] = sel_i[4] ? _1815_ : _1814_;
  assign _1816_ = sel_i[3] ? _0366_ : _0373_;
  assign _1817_ = sel_i[3] ? _0381_ : _0388_;
  assign data_o[140] = sel_i[4] ? _1817_ : _1816_;
  assign _1818_ = sel_i[3] ? _0396_ : _0403_;
  assign _1819_ = sel_i[3] ? _0411_ : _0418_;
  assign data_o[141] = sel_i[4] ? _1819_ : _1818_;
  assign _1820_ = sel_i[3] ? _0426_ : _0433_;
  assign _1821_ = sel_i[3] ? _0441_ : _0448_;
  assign data_o[142] = sel_i[4] ? _1821_ : _1820_;
  assign _1822_ = sel_i[3] ? _0456_ : _0463_;
  assign _1823_ = sel_i[3] ? _0471_ : _0478_;
  assign data_o[143] = sel_i[4] ? _1823_ : _1822_;
  assign _1824_ = sel_i[3] ? _0486_ : _0493_;
  assign _1825_ = sel_i[3] ? _0501_ : _0508_;
  assign data_o[144] = sel_i[4] ? _1825_ : _1824_;
  assign _1826_ = sel_i[3] ? _0516_ : _0523_;
  assign _1827_ = sel_i[3] ? _0531_ : _0538_;
  assign data_o[145] = sel_i[4] ? _1827_ : _1826_;
  assign _1828_ = sel_i[3] ? _0546_ : _0553_;
  assign _1829_ = sel_i[3] ? _0561_ : _0568_;
  assign data_o[146] = sel_i[4] ? _1829_ : _1828_;
  assign _1830_ = sel_i[3] ? _0576_ : _0583_;
  assign _1831_ = sel_i[3] ? _0591_ : _0598_;
  assign data_o[147] = sel_i[4] ? _1831_ : _1830_;
  assign _1832_ = sel_i[3] ? _0606_ : _0613_;
  assign _1833_ = sel_i[3] ? _0621_ : _0628_;
  assign data_o[148] = sel_i[4] ? _1833_ : _1832_;
  assign _1834_ = sel_i[3] ? _0636_ : _0643_;
  assign _1835_ = sel_i[3] ? _0651_ : _0658_;
  assign data_o[149] = sel_i[4] ? _1835_ : _1834_;
  assign _1836_ = sel_i[3] ? _0666_ : _0673_;
  assign _1837_ = sel_i[3] ? _0681_ : _0688_;
  assign data_o[150] = sel_i[4] ? _1837_ : _1836_;
  assign _1838_ = sel_i[3] ? _0696_ : _0703_;
  assign _1839_ = sel_i[3] ? _0711_ : _0718_;
  assign data_o[151] = sel_i[4] ? _1839_ : _1838_;
  assign _1840_ = sel_i[3] ? _0726_ : _0733_;
  assign _1841_ = sel_i[3] ? _0741_ : _0748_;
  assign data_o[152] = sel_i[4] ? _1841_ : _1840_;
  assign _1842_ = sel_i[3] ? _0756_ : _0763_;
  assign _1843_ = sel_i[3] ? _0771_ : _0778_;
  assign data_o[153] = sel_i[4] ? _1843_ : _1842_;
  assign _1844_ = sel_i[3] ? _0786_ : _0793_;
  assign _1845_ = sel_i[3] ? _0801_ : _0808_;
  assign data_o[154] = sel_i[4] ? _1845_ : _1844_;
  assign _1846_ = sel_i[3] ? _0816_ : _0823_;
  assign _1847_ = sel_i[3] ? _0831_ : _0838_;
  assign data_o[155] = sel_i[4] ? _1847_ : _1846_;
  assign _1848_ = sel_i[3] ? _0846_ : _0853_;
  assign _1849_ = sel_i[3] ? _0861_ : _0868_;
  assign data_o[156] = sel_i[4] ? _1849_ : _1848_;
  assign _1850_ = sel_i[3] ? _0876_ : _0883_;
  assign _1851_ = sel_i[3] ? _0891_ : _0898_;
  assign data_o[157] = sel_i[4] ? _1851_ : _1850_;
  assign _1852_ = sel_i[3] ? _0906_ : _0913_;
  assign _1853_ = sel_i[3] ? _0921_ : _0928_;
  assign data_o[158] = sel_i[4] ? _1853_ : _1852_;
  assign _1854_ = sel_i[3] ? _0936_ : _0943_;
  assign _1855_ = sel_i[3] ? _0951_ : _0958_;
  assign data_o[159] = sel_i[4] ? _1855_ : _1854_;
  assign _1856_ = sel_i[3] ? _0962_ : _0965_;
  assign _1857_ = sel_i[3] ? _0969_ : _0972_;
  assign data_o[160] = sel_i[4] ? _1857_ : _1856_;
  assign _1858_ = sel_i[3] ? _0976_ : _0979_;
  assign _1859_ = sel_i[3] ? _0983_ : _0986_;
  assign data_o[161] = sel_i[4] ? _1859_ : _1858_;
  assign _1860_ = sel_i[3] ? _0990_ : _0993_;
  assign _1861_ = sel_i[3] ? _0997_ : _1000_;
  assign data_o[162] = sel_i[4] ? _1861_ : _1860_;
  assign _1862_ = sel_i[3] ? _1004_ : _1007_;
  assign _1863_ = sel_i[3] ? _1011_ : _1014_;
  assign data_o[163] = sel_i[4] ? _1863_ : _1862_;
  assign _1864_ = sel_i[3] ? _1018_ : _1021_;
  assign _1865_ = sel_i[3] ? _1025_ : _1028_;
  assign data_o[164] = sel_i[4] ? _1865_ : _1864_;
  assign _1866_ = sel_i[3] ? _1032_ : _1035_;
  assign _1867_ = sel_i[3] ? _1039_ : _1042_;
  assign data_o[165] = sel_i[4] ? _1867_ : _1866_;
  assign _1868_ = sel_i[3] ? _1046_ : _1049_;
  assign _1869_ = sel_i[3] ? _1053_ : _1056_;
  assign data_o[166] = sel_i[4] ? _1869_ : _1868_;
  assign _1870_ = sel_i[3] ? _1060_ : _1063_;
  assign _1871_ = sel_i[3] ? _1067_ : _1070_;
  assign data_o[167] = sel_i[4] ? _1871_ : _1870_;
  assign _1872_ = sel_i[3] ? _1074_ : _1077_;
  assign _1873_ = sel_i[3] ? _1081_ : _1084_;
  assign data_o[168] = sel_i[4] ? _1873_ : _1872_;
  assign _1874_ = sel_i[3] ? _1088_ : _1091_;
  assign _1875_ = sel_i[3] ? _1095_ : _1098_;
  assign data_o[169] = sel_i[4] ? _1875_ : _1874_;
  assign _1876_ = sel_i[3] ? _1102_ : _1105_;
  assign _1877_ = sel_i[3] ? _1109_ : _1112_;
  assign data_o[170] = sel_i[4] ? _1877_ : _1876_;
  assign _1878_ = sel_i[3] ? _1116_ : _1119_;
  assign _1879_ = sel_i[3] ? _1123_ : _1126_;
  assign data_o[171] = sel_i[4] ? _1879_ : _1878_;
  assign _1880_ = sel_i[3] ? _1130_ : _1133_;
  assign _1881_ = sel_i[3] ? _1137_ : _1140_;
  assign data_o[172] = sel_i[4] ? _1881_ : _1880_;
  assign _1882_ = sel_i[3] ? _1144_ : _1147_;
  assign _1883_ = sel_i[3] ? _1151_ : _1154_;
  assign data_o[173] = sel_i[4] ? _1883_ : _1882_;
  assign _1884_ = sel_i[3] ? _1158_ : _1161_;
  assign _1885_ = sel_i[3] ? _1165_ : _1168_;
  assign data_o[174] = sel_i[4] ? _1885_ : _1884_;
  assign _1886_ = sel_i[3] ? _1172_ : _1175_;
  assign _1887_ = sel_i[3] ? _1179_ : _1182_;
  assign data_o[175] = sel_i[4] ? _1887_ : _1886_;
  assign _1888_ = sel_i[3] ? _1186_ : _1189_;
  assign _1889_ = sel_i[3] ? _1193_ : _1196_;
  assign data_o[176] = sel_i[4] ? _1889_ : _1888_;
  assign _1890_ = sel_i[3] ? _1200_ : _1203_;
  assign _1891_ = sel_i[3] ? _1207_ : _1210_;
  assign data_o[177] = sel_i[4] ? _1891_ : _1890_;
  assign _1892_ = sel_i[3] ? _1214_ : _1217_;
  assign _1893_ = sel_i[3] ? _1221_ : _1224_;
  assign data_o[178] = sel_i[4] ? _1893_ : _1892_;
  assign _1894_ = sel_i[3] ? _1228_ : _1231_;
  assign _1895_ = sel_i[3] ? _1235_ : _1238_;
  assign data_o[179] = sel_i[4] ? _1895_ : _1894_;
  assign _1896_ = sel_i[3] ? _1242_ : _1245_;
  assign _1897_ = sel_i[3] ? _1249_ : _1252_;
  assign data_o[180] = sel_i[4] ? _1897_ : _1896_;
  assign _1898_ = sel_i[3] ? _1256_ : _1259_;
  assign _1899_ = sel_i[3] ? _1263_ : _1266_;
  assign data_o[181] = sel_i[4] ? _1899_ : _1898_;
  assign _1900_ = sel_i[3] ? _1270_ : _1273_;
  assign _1901_ = sel_i[3] ? _1277_ : _1280_;
  assign data_o[182] = sel_i[4] ? _1901_ : _1900_;
  assign _1902_ = sel_i[3] ? _1284_ : _1287_;
  assign _1903_ = sel_i[3] ? _1291_ : _1294_;
  assign data_o[183] = sel_i[4] ? _1903_ : _1902_;
  assign _1904_ = sel_i[3] ? _1298_ : _1301_;
  assign _1905_ = sel_i[3] ? _1305_ : _1308_;
  assign data_o[184] = sel_i[4] ? _1905_ : _1904_;
  assign _1906_ = sel_i[3] ? _1312_ : _1315_;
  assign _1907_ = sel_i[3] ? _1319_ : _1322_;
  assign data_o[185] = sel_i[4] ? _1907_ : _1906_;
  assign _1908_ = sel_i[3] ? _1326_ : _1329_;
  assign _1909_ = sel_i[3] ? _1333_ : _1336_;
  assign data_o[186] = sel_i[4] ? _1909_ : _1908_;
  assign _1910_ = sel_i[3] ? _1340_ : _1343_;
  assign _1911_ = sel_i[3] ? _1347_ : _1350_;
  assign data_o[187] = sel_i[4] ? _1911_ : _1910_;
  assign _1912_ = sel_i[3] ? _1354_ : _1357_;
  assign _1913_ = sel_i[3] ? _1361_ : _1364_;
  assign data_o[188] = sel_i[4] ? _1913_ : _1912_;
  assign _1914_ = sel_i[3] ? _1368_ : _1371_;
  assign _1915_ = sel_i[3] ? _1375_ : _1378_;
  assign data_o[189] = sel_i[4] ? _1915_ : _1914_;
  assign _1916_ = sel_i[3] ? _1382_ : _1385_;
  assign _1917_ = sel_i[3] ? _1389_ : _1392_;
  assign data_o[190] = sel_i[4] ? _1917_ : _1916_;
  assign _1918_ = sel_i[3] ? _1396_ : _1399_;
  assign _1919_ = sel_i[3] ? _1403_ : _1406_;
  assign data_o[191] = sel_i[4] ? _1919_ : _1918_;
  assign _1920_ = sel_i[3] ? _1408_ : _1409_;
  assign _1921_ = sel_i[3] ? _1411_ : _1412_;
  assign data_o[192] = sel_i[4] ? _1921_ : _1920_;
  assign _1922_ = sel_i[3] ? _1414_ : _1415_;
  assign _1923_ = sel_i[3] ? _1417_ : _1418_;
  assign data_o[193] = sel_i[4] ? _1923_ : _1922_;
  assign _1924_ = sel_i[3] ? _1420_ : _1421_;
  assign _1925_ = sel_i[3] ? _1423_ : _1424_;
  assign data_o[194] = sel_i[4] ? _1925_ : _1924_;
  assign _1926_ = sel_i[3] ? _1426_ : _1427_;
  assign _1927_ = sel_i[3] ? _1429_ : _1430_;
  assign data_o[195] = sel_i[4] ? _1927_ : _1926_;
  assign _1928_ = sel_i[3] ? _1432_ : _1433_;
  assign _1929_ = sel_i[3] ? _1435_ : _1436_;
  assign data_o[196] = sel_i[4] ? _1929_ : _1928_;
  assign _1930_ = sel_i[3] ? _1438_ : _1439_;
  assign _1931_ = sel_i[3] ? _1441_ : _1442_;
  assign data_o[197] = sel_i[4] ? _1931_ : _1930_;
  assign _1932_ = sel_i[3] ? _1444_ : _1445_;
  assign _1933_ = sel_i[3] ? _1447_ : _1448_;
  assign data_o[198] = sel_i[4] ? _1933_ : _1932_;
  assign _1934_ = sel_i[3] ? _1450_ : _1451_;
  assign _1935_ = sel_i[3] ? _1453_ : _1454_;
  assign data_o[199] = sel_i[4] ? _1935_ : _1934_;
  assign _1936_ = sel_i[3] ? _1456_ : _1457_;
  assign _1937_ = sel_i[3] ? _1459_ : _1460_;
  assign data_o[200] = sel_i[4] ? _1937_ : _1936_;
  assign _1938_ = sel_i[3] ? _1462_ : _1463_;
  assign _1939_ = sel_i[3] ? _1465_ : _1466_;
  assign data_o[201] = sel_i[4] ? _1939_ : _1938_;
  assign _1940_ = sel_i[3] ? _1468_ : _1469_;
  assign _1941_ = sel_i[3] ? _1471_ : _1472_;
  assign data_o[202] = sel_i[4] ? _1941_ : _1940_;
  assign _1942_ = sel_i[3] ? _1474_ : _1475_;
  assign _1943_ = sel_i[3] ? _1477_ : _1478_;
  assign data_o[203] = sel_i[4] ? _1943_ : _1942_;
  assign _1944_ = sel_i[3] ? _1480_ : _1481_;
  assign _1945_ = sel_i[3] ? _1483_ : _1484_;
  assign data_o[204] = sel_i[4] ? _1945_ : _1944_;
  assign _1946_ = sel_i[3] ? _1486_ : _1487_;
  assign _1947_ = sel_i[3] ? _1489_ : _1490_;
  assign data_o[205] = sel_i[4] ? _1947_ : _1946_;
  assign _1948_ = sel_i[3] ? _1492_ : _1493_;
  assign _1949_ = sel_i[3] ? _1495_ : _1496_;
  assign data_o[206] = sel_i[4] ? _1949_ : _1948_;
  assign _1950_ = sel_i[3] ? _1498_ : _1499_;
  assign _1951_ = sel_i[3] ? _1501_ : _1502_;
  assign data_o[207] = sel_i[4] ? _1951_ : _1950_;
  assign _1952_ = sel_i[3] ? _1504_ : _1505_;
  assign _1953_ = sel_i[3] ? _1507_ : _1508_;
  assign data_o[208] = sel_i[4] ? _1953_ : _1952_;
  assign _1954_ = sel_i[3] ? _1510_ : _1511_;
  assign _1955_ = sel_i[3] ? _1513_ : _1514_;
  assign data_o[209] = sel_i[4] ? _1955_ : _1954_;
  assign _1956_ = sel_i[3] ? _1516_ : _1517_;
  assign _1957_ = sel_i[3] ? _1519_ : _1520_;
  assign data_o[210] = sel_i[4] ? _1957_ : _1956_;
  assign _1958_ = sel_i[3] ? _1522_ : _1523_;
  assign _1959_ = sel_i[3] ? _1525_ : _1526_;
  assign data_o[211] = sel_i[4] ? _1959_ : _1958_;
  assign _1960_ = sel_i[3] ? _1528_ : _1529_;
  assign _1961_ = sel_i[3] ? _1531_ : _1532_;
  assign data_o[212] = sel_i[4] ? _1961_ : _1960_;
  assign _1962_ = sel_i[3] ? _1534_ : _1535_;
  assign _1963_ = sel_i[3] ? _1537_ : _1538_;
  assign data_o[213] = sel_i[4] ? _1963_ : _1962_;
  assign _1964_ = sel_i[3] ? _1540_ : _1541_;
  assign _1965_ = sel_i[3] ? _1543_ : _1544_;
  assign data_o[214] = sel_i[4] ? _1965_ : _1964_;
  assign _1966_ = sel_i[3] ? _1546_ : _1547_;
  assign _1967_ = sel_i[3] ? _1549_ : _1550_;
  assign data_o[215] = sel_i[4] ? _1967_ : _1966_;
  assign _1968_ = sel_i[3] ? _1552_ : _1553_;
  assign _1969_ = sel_i[3] ? _1555_ : _1556_;
  assign data_o[216] = sel_i[4] ? _1969_ : _1968_;
  assign _1970_ = sel_i[3] ? _1558_ : _1559_;
  assign _1971_ = sel_i[3] ? _1561_ : _1562_;
  assign data_o[217] = sel_i[4] ? _1971_ : _1970_;
  assign _1972_ = sel_i[3] ? _1564_ : _1565_;
  assign _1973_ = sel_i[3] ? _1567_ : _1568_;
  assign data_o[218] = sel_i[4] ? _1973_ : _1972_;
  assign _1974_ = sel_i[3] ? _1570_ : _1571_;
  assign _1975_ = sel_i[3] ? _1573_ : _1574_;
  assign data_o[219] = sel_i[4] ? _1975_ : _1974_;
  assign _1976_ = sel_i[3] ? _1576_ : _1577_;
  assign _1977_ = sel_i[3] ? _1579_ : _1580_;
  assign data_o[220] = sel_i[4] ? _1977_ : _1976_;
  assign _1978_ = sel_i[3] ? _1582_ : _1583_;
  assign _1979_ = sel_i[3] ? _1585_ : _1586_;
  assign data_o[221] = sel_i[4] ? _1979_ : _1978_;
  assign _1980_ = sel_i[3] ? _1588_ : _1589_;
  assign _1981_ = sel_i[3] ? _1591_ : _1592_;
  assign data_o[222] = sel_i[4] ? _1981_ : _1980_;
  assign _1982_ = sel_i[3] ? _1594_ : _1595_;
  assign _1983_ = sel_i[3] ? _1597_ : _1598_;
  assign data_o[223] = sel_i[4] ? _1983_ : _1982_;
  assign _1984_ = sel_i[3] ? _1600_ : _1601_;
  assign _1985_ = sel_i[3] ? _1603_ : _1604_;
  assign data_o[224] = sel_i[4] ? _1985_ : _1984_;
  assign _1986_ = sel_i[3] ? _1606_ : _1607_;
  assign _1987_ = sel_i[3] ? _1609_ : _1610_;
  assign data_o[225] = sel_i[4] ? _1987_ : _1986_;
  assign _1988_ = sel_i[3] ? _1612_ : _1613_;
  assign _1989_ = sel_i[3] ? _1615_ : _1616_;
  assign data_o[226] = sel_i[4] ? _1989_ : _1988_;
  assign _1990_ = sel_i[3] ? _1618_ : _1619_;
  assign _1991_ = sel_i[3] ? _1621_ : _1622_;
  assign data_o[227] = sel_i[4] ? _1991_ : _1990_;
  assign _1992_ = sel_i[3] ? _1624_ : _1625_;
  assign _1993_ = sel_i[3] ? _1627_ : _1628_;
  assign data_o[228] = sel_i[4] ? _1993_ : _1992_;
  assign _1994_ = sel_i[3] ? _1630_ : _1631_;
  assign _1995_ = sel_i[3] ? _1633_ : _1634_;
  assign data_o[229] = sel_i[4] ? _1995_ : _1994_;
  assign _1996_ = sel_i[3] ? _1636_ : _1637_;
  assign _1997_ = sel_i[3] ? _1639_ : _1640_;
  assign data_o[230] = sel_i[4] ? _1997_ : _1996_;
  assign _1998_ = sel_i[3] ? _1642_ : _1643_;
  assign _1999_ = sel_i[3] ? _1645_ : _1646_;
  assign data_o[231] = sel_i[4] ? _1999_ : _1998_;
  assign _2000_ = sel_i[3] ? _1648_ : _1649_;
  assign _2001_ = sel_i[3] ? _1651_ : _1652_;
  assign data_o[232] = sel_i[4] ? _2001_ : _2000_;
  assign _2002_ = sel_i[3] ? _1654_ : _1655_;
  assign _2003_ = sel_i[3] ? _1657_ : _1658_;
  assign data_o[233] = sel_i[4] ? _2003_ : _2002_;
  assign _2004_ = sel_i[3] ? _1660_ : _1661_;
  assign _2005_ = sel_i[3] ? _1663_ : _1664_;
  assign data_o[234] = sel_i[4] ? _2005_ : _2004_;
  assign _2006_ = sel_i[3] ? _1666_ : _1667_;
  assign _2007_ = sel_i[3] ? _1669_ : _1670_;
  assign data_o[235] = sel_i[4] ? _2007_ : _2006_;
  assign _2008_ = sel_i[3] ? _1672_ : _1673_;
  assign _2009_ = sel_i[3] ? _1675_ : _1676_;
  assign data_o[236] = sel_i[4] ? _2009_ : _2008_;
  assign _2010_ = sel_i[3] ? _1678_ : _1679_;
  assign _2011_ = sel_i[3] ? _1681_ : _1682_;
  assign data_o[237] = sel_i[4] ? _2011_ : _2010_;
  assign _2012_ = sel_i[3] ? _1684_ : _1685_;
  assign _2013_ = sel_i[3] ? _1687_ : _1688_;
  assign data_o[238] = sel_i[4] ? _2013_ : _2012_;
  assign _2014_ = sel_i[3] ? _1690_ : _1691_;
  assign _2015_ = sel_i[3] ? _1693_ : _1694_;
  assign data_o[239] = sel_i[4] ? _2015_ : _2014_;
  assign _2016_ = sel_i[3] ? _1696_ : _1697_;
  assign _2017_ = sel_i[3] ? _1699_ : _1700_;
  assign data_o[240] = sel_i[4] ? _2017_ : _2016_;
  assign _2018_ = sel_i[3] ? _1702_ : _1703_;
  assign _2019_ = sel_i[3] ? _1705_ : _1706_;
  assign data_o[241] = sel_i[4] ? _2019_ : _2018_;
  assign _2020_ = sel_i[3] ? _1708_ : _1709_;
  assign _2021_ = sel_i[3] ? _1711_ : _1712_;
  assign data_o[242] = sel_i[4] ? _2021_ : _2020_;
  assign _2022_ = sel_i[3] ? _1714_ : _1715_;
  assign _2023_ = sel_i[3] ? _1717_ : _1718_;
  assign data_o[243] = sel_i[4] ? _2023_ : _2022_;
  assign _2024_ = sel_i[3] ? _1720_ : _1721_;
  assign _2025_ = sel_i[3] ? _1723_ : _1724_;
  assign data_o[244] = sel_i[4] ? _2025_ : _2024_;
  assign _2026_ = sel_i[3] ? _1726_ : _1727_;
  assign _2027_ = sel_i[3] ? _1729_ : _1730_;
  assign data_o[245] = sel_i[4] ? _2027_ : _2026_;
  assign _2028_ = sel_i[3] ? _1732_ : _1733_;
  assign _2029_ = sel_i[3] ? _1735_ : _1736_;
  assign data_o[246] = sel_i[4] ? _2029_ : _2028_;
  assign _2030_ = sel_i[3] ? _1738_ : _1739_;
  assign _2031_ = sel_i[3] ? _1741_ : _1742_;
  assign data_o[247] = sel_i[4] ? _2031_ : _2030_;
  assign _2032_ = sel_i[3] ? _1744_ : _1745_;
  assign _2033_ = sel_i[3] ? _1747_ : _1748_;
  assign data_o[248] = sel_i[4] ? _2033_ : _2032_;
  assign _2034_ = sel_i[3] ? _1750_ : _1751_;
  assign _2035_ = sel_i[3] ? _1753_ : _1754_;
  assign data_o[249] = sel_i[4] ? _2035_ : _2034_;
  assign _2036_ = sel_i[3] ? _1756_ : _1757_;
  assign _2037_ = sel_i[3] ? _1759_ : _1760_;
  assign data_o[250] = sel_i[4] ? _2037_ : _2036_;
  assign _2038_ = sel_i[3] ? _1762_ : _1763_;
  assign _2039_ = sel_i[3] ? _1765_ : _1766_;
  assign data_o[251] = sel_i[4] ? _2039_ : _2038_;
  assign _2040_ = sel_i[3] ? _1768_ : _1769_;
  assign _2041_ = sel_i[3] ? _1771_ : _1772_;
  assign data_o[252] = sel_i[4] ? _2041_ : _2040_;
  assign _2042_ = sel_i[3] ? _1774_ : _1775_;
  assign _2043_ = sel_i[3] ? _1777_ : _1778_;
  assign data_o[253] = sel_i[4] ? _2043_ : _2042_;
  assign _2044_ = sel_i[3] ? _1780_ : _1781_;
  assign _2045_ = sel_i[3] ? _1783_ : _1784_;
  assign data_o[254] = sel_i[4] ? _2045_ : _2044_;
  assign _2046_ = sel_i[3] ? _1786_ : _1787_;
  assign _2047_ = sel_i[3] ? _1789_ : _1790_;
  assign data_o[255] = sel_i[4] ? _2047_ : _2046_;
  assign data_o[256] = sel_i[4] ? _0014_ : _0029_;
  assign data_o[257] = sel_i[4] ? _0044_ : _0059_;
  assign data_o[258] = sel_i[4] ? _0074_ : _0089_;
  assign data_o[259] = sel_i[4] ? _0104_ : _0119_;
  assign data_o[260] = sel_i[4] ? _0134_ : _0149_;
  assign data_o[261] = sel_i[4] ? _0164_ : _0179_;
  assign data_o[262] = sel_i[4] ? _0194_ : _0209_;
  assign data_o[263] = sel_i[4] ? _0224_ : _0239_;
  assign data_o[264] = sel_i[4] ? _0254_ : _0269_;
  assign data_o[265] = sel_i[4] ? _0284_ : _0299_;
  assign data_o[266] = sel_i[4] ? _0314_ : _0329_;
  assign data_o[267] = sel_i[4] ? _0344_ : _0359_;
  assign data_o[268] = sel_i[4] ? _0374_ : _0389_;
  assign data_o[269] = sel_i[4] ? _0404_ : _0419_;
  assign data_o[270] = sel_i[4] ? _0434_ : _0449_;
  assign data_o[271] = sel_i[4] ? _0464_ : _0479_;
  assign data_o[272] = sel_i[4] ? _0494_ : _0509_;
  assign data_o[273] = sel_i[4] ? _0524_ : _0539_;
  assign data_o[274] = sel_i[4] ? _0554_ : _0569_;
  assign data_o[275] = sel_i[4] ? _0584_ : _0599_;
  assign data_o[276] = sel_i[4] ? _0614_ : _0629_;
  assign data_o[277] = sel_i[4] ? _0644_ : _0659_;
  assign data_o[278] = sel_i[4] ? _0674_ : _0689_;
  assign data_o[279] = sel_i[4] ? _0704_ : _0719_;
  assign data_o[280] = sel_i[4] ? _0734_ : _0749_;
  assign data_o[281] = sel_i[4] ? _0764_ : _0779_;
  assign data_o[282] = sel_i[4] ? _0794_ : _0809_;
  assign data_o[283] = sel_i[4] ? _0824_ : _0839_;
  assign data_o[284] = sel_i[4] ? _0854_ : _0869_;
  assign data_o[285] = sel_i[4] ? _0884_ : _0899_;
  assign data_o[286] = sel_i[4] ? _0914_ : _0929_;
  assign data_o[287] = sel_i[4] ? _0944_ : _0959_;
  assign data_o[288] = sel_i[4] ? _0966_ : _0973_;
  assign data_o[289] = sel_i[4] ? _0980_ : _0987_;
  assign data_o[290] = sel_i[4] ? _0994_ : _1001_;
  assign data_o[291] = sel_i[4] ? _1008_ : _1015_;
  assign data_o[292] = sel_i[4] ? _1022_ : _1029_;
  assign data_o[293] = sel_i[4] ? _1036_ : _1043_;
  assign data_o[294] = sel_i[4] ? _1050_ : _1057_;
  assign data_o[295] = sel_i[4] ? _1064_ : _1071_;
  assign data_o[296] = sel_i[4] ? _1078_ : _1085_;
  assign data_o[297] = sel_i[4] ? _1092_ : _1099_;
  assign data_o[298] = sel_i[4] ? _1106_ : _1113_;
  assign data_o[299] = sel_i[4] ? _1120_ : _1127_;
  assign data_o[300] = sel_i[4] ? _1134_ : _1141_;
  assign data_o[301] = sel_i[4] ? _1148_ : _1155_;
  assign data_o[302] = sel_i[4] ? _1162_ : _1169_;
  assign data_o[303] = sel_i[4] ? _1176_ : _1183_;
  assign data_o[304] = sel_i[4] ? _1190_ : _1197_;
  assign data_o[305] = sel_i[4] ? _1204_ : _1211_;
  assign data_o[306] = sel_i[4] ? _1218_ : _1225_;
  assign data_o[307] = sel_i[4] ? _1232_ : _1239_;
  assign data_o[308] = sel_i[4] ? _1246_ : _1253_;
  assign data_o[309] = sel_i[4] ? _1260_ : _1267_;
  assign data_o[310] = sel_i[4] ? _1274_ : _1281_;
  assign data_o[311] = sel_i[4] ? _1288_ : _1295_;
  assign data_o[312] = sel_i[4] ? _1302_ : _1309_;
  assign data_o[313] = sel_i[4] ? _1316_ : _1323_;
  assign data_o[314] = sel_i[4] ? _1330_ : _1337_;
  assign data_o[315] = sel_i[4] ? _1344_ : _1351_;
  assign data_o[316] = sel_i[4] ? _1358_ : _1365_;
  assign data_o[317] = sel_i[4] ? _1372_ : _1379_;
  assign data_o[318] = sel_i[4] ? _1386_ : _1393_;
  assign data_o[319] = sel_i[4] ? _1400_ : _1407_;
  assign data_o[320] = sel_i[4] ? _1410_ : _1413_;
  assign data_o[321] = sel_i[4] ? _1416_ : _1419_;
  assign data_o[322] = sel_i[4] ? _1422_ : _1425_;
  assign data_o[323] = sel_i[4] ? _1428_ : _1431_;
  assign data_o[324] = sel_i[4] ? _1434_ : _1437_;
  assign data_o[325] = sel_i[4] ? _1440_ : _1443_;
  assign data_o[326] = sel_i[4] ? _1446_ : _1449_;
  assign data_o[327] = sel_i[4] ? _1452_ : _1455_;
  assign data_o[328] = sel_i[4] ? _1458_ : _1461_;
  assign data_o[329] = sel_i[4] ? _1464_ : _1467_;
  assign data_o[330] = sel_i[4] ? _1470_ : _1473_;
  assign data_o[331] = sel_i[4] ? _1476_ : _1479_;
  assign data_o[332] = sel_i[4] ? _1482_ : _1485_;
  assign data_o[333] = sel_i[4] ? _1488_ : _1491_;
  assign data_o[334] = sel_i[4] ? _1494_ : _1497_;
  assign data_o[335] = sel_i[4] ? _1500_ : _1503_;
  assign data_o[336] = sel_i[4] ? _1506_ : _1509_;
  assign data_o[337] = sel_i[4] ? _1512_ : _1515_;
  assign data_o[338] = sel_i[4] ? _1518_ : _1521_;
  assign data_o[339] = sel_i[4] ? _1524_ : _1527_;
  assign data_o[340] = sel_i[4] ? _1530_ : _1533_;
  assign data_o[341] = sel_i[4] ? _1536_ : _1539_;
  assign data_o[342] = sel_i[4] ? _1542_ : _1545_;
  assign data_o[343] = sel_i[4] ? _1548_ : _1551_;
  assign data_o[344] = sel_i[4] ? _1554_ : _1557_;
  assign data_o[345] = sel_i[4] ? _1560_ : _1563_;
  assign data_o[346] = sel_i[4] ? _1566_ : _1569_;
  assign data_o[347] = sel_i[4] ? _1572_ : _1575_;
  assign data_o[348] = sel_i[4] ? _1578_ : _1581_;
  assign data_o[349] = sel_i[4] ? _1584_ : _1587_;
  assign data_o[350] = sel_i[4] ? _1590_ : _1593_;
  assign data_o[351] = sel_i[4] ? _1596_ : _1599_;
  assign data_o[352] = sel_i[4] ? _1602_ : _1605_;
  assign data_o[353] = sel_i[4] ? _1608_ : _1611_;
  assign data_o[354] = sel_i[4] ? _1614_ : _1617_;
  assign data_o[355] = sel_i[4] ? _1620_ : _1623_;
  assign data_o[356] = sel_i[4] ? _1626_ : _1629_;
  assign data_o[357] = sel_i[4] ? _1632_ : _1635_;
  assign data_o[358] = sel_i[4] ? _1638_ : _1641_;
  assign data_o[359] = sel_i[4] ? _1644_ : _1647_;
  assign data_o[360] = sel_i[4] ? _1650_ : _1653_;
  assign data_o[361] = sel_i[4] ? _1656_ : _1659_;
  assign data_o[362] = sel_i[4] ? _1662_ : _1665_;
  assign data_o[363] = sel_i[4] ? _1668_ : _1671_;
  assign data_o[364] = sel_i[4] ? _1674_ : _1677_;
  assign data_o[365] = sel_i[4] ? _1680_ : _1683_;
  assign data_o[366] = sel_i[4] ? _1686_ : _1689_;
  assign data_o[367] = sel_i[4] ? _1692_ : _1695_;
  assign data_o[368] = sel_i[4] ? _1698_ : _1701_;
  assign data_o[369] = sel_i[4] ? _1704_ : _1707_;
  assign data_o[370] = sel_i[4] ? _1710_ : _1713_;
  assign data_o[371] = sel_i[4] ? _1716_ : _1719_;
  assign data_o[372] = sel_i[4] ? _1722_ : _1725_;
  assign data_o[373] = sel_i[4] ? _1728_ : _1731_;
  assign data_o[374] = sel_i[4] ? _1734_ : _1737_;
  assign data_o[375] = sel_i[4] ? _1740_ : _1743_;
  assign data_o[376] = sel_i[4] ? _1746_ : _1749_;
  assign data_o[377] = sel_i[4] ? _1752_ : _1755_;
  assign data_o[378] = sel_i[4] ? _1758_ : _1761_;
  assign data_o[379] = sel_i[4] ? _1764_ : _1767_;
  assign data_o[380] = sel_i[4] ? _1770_ : _1773_;
  assign data_o[381] = sel_i[4] ? _1776_ : _1779_;
  assign data_o[382] = sel_i[4] ? _1782_ : _1785_;
  assign data_o[383] = sel_i[4] ? _1788_ : _1791_;
  assign data_o[384] = sel_i[4] ? _1792_ : _1793_;
  assign data_o[385] = sel_i[4] ? _1794_ : _1795_;
  assign data_o[386] = sel_i[4] ? _1796_ : _1797_;
  assign data_o[387] = sel_i[4] ? _1798_ : _1799_;
  assign data_o[388] = sel_i[4] ? _1800_ : _1801_;
  assign data_o[389] = sel_i[4] ? _1802_ : _1803_;
  assign data_o[390] = sel_i[4] ? _1804_ : _1805_;
  assign data_o[391] = sel_i[4] ? _1806_ : _1807_;
  assign data_o[392] = sel_i[4] ? _1808_ : _1809_;
  assign data_o[393] = sel_i[4] ? _1810_ : _1811_;
  assign data_o[394] = sel_i[4] ? _1812_ : _1813_;
  assign data_o[395] = sel_i[4] ? _1814_ : _1815_;
  assign data_o[396] = sel_i[4] ? _1816_ : _1817_;
  assign data_o[397] = sel_i[4] ? _1818_ : _1819_;
  assign data_o[398] = sel_i[4] ? _1820_ : _1821_;
  assign data_o[399] = sel_i[4] ? _1822_ : _1823_;
  assign data_o[400] = sel_i[4] ? _1824_ : _1825_;
  assign data_o[401] = sel_i[4] ? _1826_ : _1827_;
  assign data_o[402] = sel_i[4] ? _1828_ : _1829_;
  assign data_o[403] = sel_i[4] ? _1830_ : _1831_;
  assign data_o[404] = sel_i[4] ? _1832_ : _1833_;
  assign data_o[405] = sel_i[4] ? _1834_ : _1835_;
  assign data_o[406] = sel_i[4] ? _1836_ : _1837_;
  assign data_o[407] = sel_i[4] ? _1838_ : _1839_;
  assign data_o[408] = sel_i[4] ? _1840_ : _1841_;
  assign data_o[409] = sel_i[4] ? _1842_ : _1843_;
  assign data_o[410] = sel_i[4] ? _1844_ : _1845_;
  assign data_o[411] = sel_i[4] ? _1846_ : _1847_;
  assign data_o[412] = sel_i[4] ? _1848_ : _1849_;
  assign data_o[413] = sel_i[4] ? _1850_ : _1851_;
  assign data_o[414] = sel_i[4] ? _1852_ : _1853_;
  assign data_o[415] = sel_i[4] ? _1854_ : _1855_;
  assign data_o[416] = sel_i[4] ? _1856_ : _1857_;
  assign data_o[417] = sel_i[4] ? _1858_ : _1859_;
  assign data_o[418] = sel_i[4] ? _1860_ : _1861_;
  assign data_o[419] = sel_i[4] ? _1862_ : _1863_;
  assign data_o[420] = sel_i[4] ? _1864_ : _1865_;
  assign data_o[421] = sel_i[4] ? _1866_ : _1867_;
  assign data_o[422] = sel_i[4] ? _1868_ : _1869_;
  assign data_o[423] = sel_i[4] ? _1870_ : _1871_;
  assign data_o[424] = sel_i[4] ? _1872_ : _1873_;
  assign data_o[425] = sel_i[4] ? _1874_ : _1875_;
  assign data_o[426] = sel_i[4] ? _1876_ : _1877_;
  assign data_o[427] = sel_i[4] ? _1878_ : _1879_;
  assign data_o[428] = sel_i[4] ? _1880_ : _1881_;
  assign data_o[429] = sel_i[4] ? _1882_ : _1883_;
  assign data_o[430] = sel_i[4] ? _1884_ : _1885_;
  assign data_o[431] = sel_i[4] ? _1886_ : _1887_;
  assign data_o[432] = sel_i[4] ? _1888_ : _1889_;
  assign data_o[433] = sel_i[4] ? _1890_ : _1891_;
  assign data_o[434] = sel_i[4] ? _1892_ : _1893_;
  assign data_o[435] = sel_i[4] ? _1894_ : _1895_;
  assign data_o[436] = sel_i[4] ? _1896_ : _1897_;
  assign data_o[437] = sel_i[4] ? _1898_ : _1899_;
  assign data_o[438] = sel_i[4] ? _1900_ : _1901_;
  assign data_o[439] = sel_i[4] ? _1902_ : _1903_;
  assign data_o[440] = sel_i[4] ? _1904_ : _1905_;
  assign data_o[441] = sel_i[4] ? _1906_ : _1907_;
  assign data_o[442] = sel_i[4] ? _1908_ : _1909_;
  assign data_o[443] = sel_i[4] ? _1910_ : _1911_;
  assign data_o[444] = sel_i[4] ? _1912_ : _1913_;
  assign data_o[445] = sel_i[4] ? _1914_ : _1915_;
  assign data_o[446] = sel_i[4] ? _1916_ : _1917_;
  assign data_o[447] = sel_i[4] ? _1918_ : _1919_;
  assign data_o[448] = sel_i[4] ? _1920_ : _1921_;
  assign data_o[449] = sel_i[4] ? _1922_ : _1923_;
  assign data_o[450] = sel_i[4] ? _1924_ : _1925_;
  assign data_o[451] = sel_i[4] ? _1926_ : _1927_;
  assign data_o[452] = sel_i[4] ? _1928_ : _1929_;
  assign data_o[453] = sel_i[4] ? _1930_ : _1931_;
  assign data_o[454] = sel_i[4] ? _1932_ : _1933_;
  assign data_o[455] = sel_i[4] ? _1934_ : _1935_;
  assign data_o[456] = sel_i[4] ? _1936_ : _1937_;
  assign data_o[457] = sel_i[4] ? _1938_ : _1939_;
  assign data_o[458] = sel_i[4] ? _1940_ : _1941_;
  assign data_o[459] = sel_i[4] ? _1942_ : _1943_;
  assign data_o[460] = sel_i[4] ? _1944_ : _1945_;
  assign data_o[461] = sel_i[4] ? _1946_ : _1947_;
  assign data_o[462] = sel_i[4] ? _1948_ : _1949_;
  assign data_o[463] = sel_i[4] ? _1950_ : _1951_;
  assign data_o[464] = sel_i[4] ? _1952_ : _1953_;
  assign data_o[465] = sel_i[4] ? _1954_ : _1955_;
  assign data_o[466] = sel_i[4] ? _1956_ : _1957_;
  assign data_o[467] = sel_i[4] ? _1958_ : _1959_;
  assign data_o[468] = sel_i[4] ? _1960_ : _1961_;
  assign data_o[469] = sel_i[4] ? _1962_ : _1963_;
  assign data_o[470] = sel_i[4] ? _1964_ : _1965_;
  assign data_o[471] = sel_i[4] ? _1966_ : _1967_;
  assign data_o[472] = sel_i[4] ? _1968_ : _1969_;
  assign data_o[473] = sel_i[4] ? _1970_ : _1971_;
  assign data_o[474] = sel_i[4] ? _1972_ : _1973_;
  assign data_o[475] = sel_i[4] ? _1974_ : _1975_;
  assign data_o[476] = sel_i[4] ? _1976_ : _1977_;
  assign data_o[477] = sel_i[4] ? _1978_ : _1979_;
  assign data_o[478] = sel_i[4] ? _1980_ : _1981_;
  assign data_o[479] = sel_i[4] ? _1982_ : _1983_;
  assign data_o[480] = sel_i[4] ? _1984_ : _1985_;
  assign data_o[481] = sel_i[4] ? _1986_ : _1987_;
  assign data_o[482] = sel_i[4] ? _1988_ : _1989_;
  assign data_o[483] = sel_i[4] ? _1990_ : _1991_;
  assign data_o[484] = sel_i[4] ? _1992_ : _1993_;
  assign data_o[485] = sel_i[4] ? _1994_ : _1995_;
  assign data_o[486] = sel_i[4] ? _1996_ : _1997_;
  assign data_o[487] = sel_i[4] ? _1998_ : _1999_;
  assign data_o[488] = sel_i[4] ? _2000_ : _2001_;
  assign data_o[489] = sel_i[4] ? _2002_ : _2003_;
  assign data_o[490] = sel_i[4] ? _2004_ : _2005_;
  assign data_o[491] = sel_i[4] ? _2006_ : _2007_;
  assign data_o[492] = sel_i[4] ? _2008_ : _2009_;
  assign data_o[493] = sel_i[4] ? _2010_ : _2011_;
  assign data_o[494] = sel_i[4] ? _2012_ : _2013_;
  assign data_o[495] = sel_i[4] ? _2014_ : _2015_;
  assign data_o[496] = sel_i[4] ? _2016_ : _2017_;
  assign data_o[497] = sel_i[4] ? _2018_ : _2019_;
  assign data_o[498] = sel_i[4] ? _2020_ : _2021_;
  assign data_o[499] = sel_i[4] ? _2022_ : _2023_;
  assign data_o[500] = sel_i[4] ? _2024_ : _2025_;
  assign data_o[501] = sel_i[4] ? _2026_ : _2027_;
  assign data_o[502] = sel_i[4] ? _2028_ : _2029_;
  assign data_o[503] = sel_i[4] ? _2030_ : _2031_;
  assign data_o[504] = sel_i[4] ? _2032_ : _2033_;
  assign data_o[505] = sel_i[4] ? _2034_ : _2035_;
  assign data_o[506] = sel_i[4] ? _2036_ : _2037_;
  assign data_o[507] = sel_i[4] ? _2038_ : _2039_;
  assign data_o[508] = sel_i[4] ? _2040_ : _2041_;
  assign data_o[509] = sel_i[4] ? _2042_ : _2043_;
  assign data_o[510] = sel_i[4] ? _2044_ : _2045_;
  assign data_o[511] = sel_i[4] ? _2046_ : _2047_;
  assign data_stage = { data_o, \mux_stage[3].mux_swap[1].swap_inst.data_o , \mux_stage[3].mux_swap[0].swap_inst.data_o , \mux_stage[2].mux_swap[3].swap_inst.data_o , \mux_stage[2].mux_swap[2].swap_inst.data_o , \mux_stage[2].mux_swap[1].swap_inst.data_o , \mux_stage[2].mux_swap[0].swap_inst.data_o , \mux_stage[1].mux_swap[7].swap_inst.data_o , \mux_stage[1].mux_swap[6].swap_inst.data_o , \mux_stage[1].mux_swap[5].swap_inst.data_o , \mux_stage[1].mux_swap[4].swap_inst.data_o , \mux_stage[1].mux_swap[3].swap_inst.data_o , \mux_stage[1].mux_swap[2].swap_inst.data_o , \mux_stage[1].mux_swap[1].swap_inst.data_o , \mux_stage[1].mux_swap[0].swap_inst.data_o , \mux_stage[0].mux_swap[15].swap_inst.data_o , \mux_stage[0].mux_swap[14].swap_inst.data_o , \mux_stage[0].mux_swap[13].swap_inst.data_o , \mux_stage[0].mux_swap[12].swap_inst.data_o , \mux_stage[0].mux_swap[11].swap_inst.data_o , \mux_stage[0].mux_swap[10].swap_inst.data_o , \mux_stage[0].mux_swap[9].swap_inst.data_o , \mux_stage[0].mux_swap[8].swap_inst.data_o , \mux_stage[0].mux_swap[7].swap_inst.data_o , \mux_stage[0].mux_swap[6].swap_inst.data_o , \mux_stage[0].mux_swap[5].swap_inst.data_o , \mux_stage[0].mux_swap[4].swap_inst.data_o , \mux_stage[0].mux_swap[3].swap_inst.data_o , \mux_stage[0].mux_swap[2].swap_inst.data_o , \mux_stage[0].mux_swap[1].swap_inst.data_o , \mux_stage[0].mux_swap[0].swap_inst.data_o , data_i };
  assign \mux_stage[0].mux_swap[0].swap_inst.data_i  = data_i[31:0];
  assign \mux_stage[0].mux_swap[0].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[10].swap_inst.data_i  = data_i[351:320];
  assign \mux_stage[0].mux_swap[10].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[11].swap_inst.data_i  = data_i[383:352];
  assign \mux_stage[0].mux_swap[11].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[12].swap_inst.data_i  = data_i[415:384];
  assign \mux_stage[0].mux_swap[12].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[13].swap_inst.data_i  = data_i[447:416];
  assign \mux_stage[0].mux_swap[13].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[14].swap_inst.data_i  = data_i[479:448];
  assign \mux_stage[0].mux_swap[14].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[15].swap_inst.data_i  = data_i[511:480];
  assign \mux_stage[0].mux_swap[15].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[1].swap_inst.data_i  = data_i[63:32];
  assign \mux_stage[0].mux_swap[1].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[2].swap_inst.data_i  = data_i[95:64];
  assign \mux_stage[0].mux_swap[2].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[3].swap_inst.data_i  = data_i[127:96];
  assign \mux_stage[0].mux_swap[3].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[4].swap_inst.data_i  = data_i[159:128];
  assign \mux_stage[0].mux_swap[4].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[5].swap_inst.data_i  = data_i[191:160];
  assign \mux_stage[0].mux_swap[5].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[6].swap_inst.data_i  = data_i[223:192];
  assign \mux_stage[0].mux_swap[6].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[7].swap_inst.data_i  = data_i[255:224];
  assign \mux_stage[0].mux_swap[7].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[8].swap_inst.data_i  = data_i[287:256];
  assign \mux_stage[0].mux_swap[8].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[0].mux_swap[9].swap_inst.data_i  = data_i[319:288];
  assign \mux_stage[0].mux_swap[9].swap_inst.swap_i  = sel_i[0];
  assign \mux_stage[1].mux_swap[0].swap_inst.data_i  = { \mux_stage[0].mux_swap[1].swap_inst.data_o , \mux_stage[0].mux_swap[0].swap_inst.data_o  };
  assign \mux_stage[1].mux_swap[0].swap_inst.swap_i  = sel_i[1];
  assign \mux_stage[1].mux_swap[1].swap_inst.data_i  = { \mux_stage[0].mux_swap[3].swap_inst.data_o , \mux_stage[0].mux_swap[2].swap_inst.data_o  };
  assign \mux_stage[1].mux_swap[1].swap_inst.swap_i  = sel_i[1];
  assign \mux_stage[1].mux_swap[2].swap_inst.data_i  = { \mux_stage[0].mux_swap[5].swap_inst.data_o , \mux_stage[0].mux_swap[4].swap_inst.data_o  };
  assign \mux_stage[1].mux_swap[2].swap_inst.swap_i  = sel_i[1];
  assign \mux_stage[1].mux_swap[3].swap_inst.data_i  = { \mux_stage[0].mux_swap[7].swap_inst.data_o , \mux_stage[0].mux_swap[6].swap_inst.data_o  };
  assign \mux_stage[1].mux_swap[3].swap_inst.swap_i  = sel_i[1];
  assign \mux_stage[1].mux_swap[4].swap_inst.data_i  = { \mux_stage[0].mux_swap[9].swap_inst.data_o , \mux_stage[0].mux_swap[8].swap_inst.data_o  };
  assign \mux_stage[1].mux_swap[4].swap_inst.swap_i  = sel_i[1];
  assign \mux_stage[1].mux_swap[5].swap_inst.data_i  = { \mux_stage[0].mux_swap[11].swap_inst.data_o , \mux_stage[0].mux_swap[10].swap_inst.data_o  };
  assign \mux_stage[1].mux_swap[5].swap_inst.swap_i  = sel_i[1];
  assign \mux_stage[1].mux_swap[6].swap_inst.data_i  = { \mux_stage[0].mux_swap[13].swap_inst.data_o , \mux_stage[0].mux_swap[12].swap_inst.data_o  };
  assign \mux_stage[1].mux_swap[6].swap_inst.swap_i  = sel_i[1];
  assign \mux_stage[1].mux_swap[7].swap_inst.data_i  = { \mux_stage[0].mux_swap[15].swap_inst.data_o , \mux_stage[0].mux_swap[14].swap_inst.data_o  };
  assign \mux_stage[1].mux_swap[7].swap_inst.swap_i  = sel_i[1];
  assign \mux_stage[2].mux_swap[0].swap_inst.data_i  = { \mux_stage[1].mux_swap[1].swap_inst.data_o , \mux_stage[1].mux_swap[0].swap_inst.data_o  };
  assign \mux_stage[2].mux_swap[0].swap_inst.swap_i  = sel_i[2];
  assign \mux_stage[2].mux_swap[1].swap_inst.data_i  = { \mux_stage[1].mux_swap[3].swap_inst.data_o , \mux_stage[1].mux_swap[2].swap_inst.data_o  };
  assign \mux_stage[2].mux_swap[1].swap_inst.swap_i  = sel_i[2];
  assign \mux_stage[2].mux_swap[2].swap_inst.data_i  = { \mux_stage[1].mux_swap[5].swap_inst.data_o , \mux_stage[1].mux_swap[4].swap_inst.data_o  };
  assign \mux_stage[2].mux_swap[2].swap_inst.swap_i  = sel_i[2];
  assign \mux_stage[2].mux_swap[3].swap_inst.data_i  = { \mux_stage[1].mux_swap[7].swap_inst.data_o , \mux_stage[1].mux_swap[6].swap_inst.data_o  };
  assign \mux_stage[2].mux_swap[3].swap_inst.swap_i  = sel_i[2];
  assign \mux_stage[3].mux_swap[0].swap_inst.data_i  = { \mux_stage[2].mux_swap[1].swap_inst.data_o , \mux_stage[2].mux_swap[0].swap_inst.data_o  };
  assign \mux_stage[3].mux_swap[0].swap_inst.swap_i  = sel_i[3];
  assign \mux_stage[3].mux_swap[1].swap_inst.data_i  = { \mux_stage[2].mux_swap[3].swap_inst.data_o , \mux_stage[2].mux_swap[2].swap_inst.data_o  };
  assign \mux_stage[3].mux_swap[1].swap_inst.swap_i  = sel_i[3];
  assign \mux_stage[4].mux_swap[0].swap_inst.data_i  = { \mux_stage[3].mux_swap[1].swap_inst.data_o , \mux_stage[3].mux_swap[0].swap_inst.data_o  };
  assign \mux_stage[4].mux_swap[0].swap_inst.data_o  = data_o;
  assign \mux_stage[4].mux_swap[0].swap_inst.swap_i  = sel_i[4];
endmodule
