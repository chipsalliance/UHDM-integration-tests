

module dut;
   undefined undef(.in('0));
endmodule
