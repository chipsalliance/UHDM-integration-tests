module bsg_fifo_tracker(clk_i, reset_i, enq_i, deq_i, wptr_r_o, rptr_r_o, rptr_n_o, full_o, empty_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  input clk_i;
  wire clk_i;
  input deq_i;
  wire deq_i;
  reg deq_r;
  wire empty;
  output empty_o;
  wire empty_o;
  input enq_i;
  wire enq_i;
  reg enq_r;
  wire full;
  output full_o;
  wire full_o;
  input reset_i;
  wire reset_i;
  wire \rptr.add_i ;
  wire \rptr.clk ;
  wire [5:0] \rptr.n_o ;
  wire [5:0] \rptr.o ;
  wire [5:0] \rptr.ptr_n ;
  reg [5:0] \rptr.ptr_r ;
  wire \rptr.reset_i ;
  wire [5:0] rptr_n;
  output [5:0] rptr_n_o;
  wire [5:0] rptr_n_o;
  wire [5:0] rptr_r;
  output [5:0] rptr_r_o;
  wire [5:0] rptr_r_o;
  wire \wptr.add_i ;
  wire \wptr.clk ;
  wire [5:0] \wptr.genblk1.genblk1.ptr_r_p1 ;
  wire [5:0] \wptr.o ;
  reg [5:0] \wptr.ptr_r ;
  wire \wptr.reset_i ;
  wire [5:0] wptr_r;
  output [5:0] wptr_r_o;
  wire [5:0] wptr_r_o;
  assign rptr_n_o[0] = deq_i ^ \rptr.ptr_r [0];
  assign _00_ = \rptr.ptr_r [1] ^ \rptr.ptr_r [0];
  assign rptr_n_o[1] = deq_i ? _00_ : \rptr.ptr_r [1];
  assign _01_ = ~(\rptr.ptr_r [1] & \rptr.ptr_r [0]);
  assign _02_ = ~(_01_ ^ \rptr.ptr_r [2]);
  assign rptr_n_o[2] = deq_i ? _02_ : \rptr.ptr_r [2];
  assign _03_ = \rptr.ptr_r [2] & ~(_01_);
  assign _04_ = _03_ ^ \rptr.ptr_r [3];
  assign rptr_n_o[3] = deq_i ? _04_ : \rptr.ptr_r [3];
  assign _05_ = ~(\rptr.ptr_r [3] & \rptr.ptr_r [2]);
  assign _06_ = _05_ | _01_;
  assign _07_ = ~(_06_ ^ \rptr.ptr_r [4]);
  assign rptr_n_o[4] = deq_i ? _07_ : \rptr.ptr_r [4];
  assign _08_ = \rptr.ptr_r [4] & ~(_06_);
  assign _09_ = _08_ ^ \rptr.ptr_r [5];
  assign rptr_n_o[5] = deq_i ? _09_ : \rptr.ptr_r [5];
  assign \wptr.genblk1.genblk1.ptr_r_p1 [0] = ~\wptr.ptr_r [0];
  assign _10_ = \wptr.ptr_r [0] ^ \rptr.ptr_r [0];
  assign _11_ = \wptr.ptr_r [1] ^ \rptr.ptr_r [1];
  assign _12_ = _11_ | _10_;
  assign _13_ = \wptr.ptr_r [2] ^ \rptr.ptr_r [2];
  assign _14_ = \wptr.ptr_r [3] ^ \rptr.ptr_r [3];
  assign _15_ = _14_ | _13_;
  assign _16_ = _15_ | _12_;
  assign _17_ = \wptr.ptr_r [4] ^ \rptr.ptr_r [4];
  assign _18_ = \wptr.ptr_r [5] ^ \rptr.ptr_r [5];
  assign _19_ = _18_ | _17_;
  assign _20_ = _19_ | _16_;
  assign empty_o = deq_r & ~(_20_);
  assign full_o = enq_r & ~(_20_);
  assign _26_ = enq_i | deq_i;
  assign \wptr.genblk1.genblk1.ptr_r_p1 [1] = \wptr.ptr_r [1] ^ \wptr.ptr_r [0];
  assign _21_ = ~(\wptr.ptr_r [1] & \wptr.ptr_r [0]);
  assign \wptr.genblk1.genblk1.ptr_r_p1 [2] = ~(_21_ ^ \wptr.ptr_r [2]);
  assign _22_ = \wptr.ptr_r [2] & ~(_21_);
  assign \wptr.genblk1.genblk1.ptr_r_p1 [3] = _22_ ^ \wptr.ptr_r [3];
  assign _23_ = ~(\wptr.ptr_r [3] & \wptr.ptr_r [2]);
  assign _24_ = _23_ | _21_;
  assign \wptr.genblk1.genblk1.ptr_r_p1 [4] = ~(_24_ ^ \wptr.ptr_r [4]);
  assign _25_ = \wptr.ptr_r [4] & ~(_24_);
  assign \wptr.genblk1.genblk1.ptr_r_p1 [5] = _25_ ^ \wptr.ptr_r [5];
  always @(posedge clk_i)
    if (reset_i) enq_r <= 1'h0;
    else if (_26_) enq_r <= enq_i;
  always @(posedge clk_i)
    if (reset_i) deq_r <= 1'h1;
    else if (_26_) deq_r <= deq_i;
  always @(posedge clk_i)
    if (reset_i) \rptr.ptr_r [0] <= 1'h0;
    else \rptr.ptr_r [0] <= rptr_n_o[0];
  always @(posedge clk_i)
    if (reset_i) \rptr.ptr_r [1] <= 1'h0;
    else \rptr.ptr_r [1] <= rptr_n_o[1];
  always @(posedge clk_i)
    if (reset_i) \rptr.ptr_r [2] <= 1'h0;
    else \rptr.ptr_r [2] <= rptr_n_o[2];
  always @(posedge clk_i)
    if (reset_i) \rptr.ptr_r [3] <= 1'h0;
    else \rptr.ptr_r [3] <= rptr_n_o[3];
  always @(posedge clk_i)
    if (reset_i) \rptr.ptr_r [4] <= 1'h0;
    else \rptr.ptr_r [4] <= rptr_n_o[4];
  always @(posedge clk_i)
    if (reset_i) \rptr.ptr_r [5] <= 1'h0;
    else \rptr.ptr_r [5] <= rptr_n_o[5];
  always @(posedge clk_i)
    if (reset_i) \wptr.ptr_r [0] <= 1'h0;
    else if (enq_i) \wptr.ptr_r [0] <= \wptr.genblk1.genblk1.ptr_r_p1 [0];
  always @(posedge clk_i)
    if (reset_i) \wptr.ptr_r [1] <= 1'h0;
    else if (enq_i) \wptr.ptr_r [1] <= \wptr.genblk1.genblk1.ptr_r_p1 [1];
  always @(posedge clk_i)
    if (reset_i) \wptr.ptr_r [2] <= 1'h0;
    else if (enq_i) \wptr.ptr_r [2] <= \wptr.genblk1.genblk1.ptr_r_p1 [2];
  always @(posedge clk_i)
    if (reset_i) \wptr.ptr_r [3] <= 1'h0;
    else if (enq_i) \wptr.ptr_r [3] <= \wptr.genblk1.genblk1.ptr_r_p1 [3];
  always @(posedge clk_i)
    if (reset_i) \wptr.ptr_r [4] <= 1'h0;
    else if (enq_i) \wptr.ptr_r [4] <= \wptr.genblk1.genblk1.ptr_r_p1 [4];
  always @(posedge clk_i)
    if (reset_i) \wptr.ptr_r [5] <= 1'h0;
    else if (enq_i) \wptr.ptr_r [5] <= \wptr.genblk1.genblk1.ptr_r_p1 [5];
  assign empty = empty_o;
  assign full = full_o;
  assign \rptr.add_i  = deq_i;
  assign \rptr.clk  = clk_i;
  assign \rptr.n_o  = rptr_n_o;
  assign \rptr.o  = \rptr.ptr_r ;
  assign \rptr.ptr_n  = rptr_n_o;
  assign \rptr.reset_i  = reset_i;
  assign rptr_n = rptr_n_o;
  assign rptr_r = \rptr.ptr_r ;
  assign rptr_r_o = \rptr.ptr_r ;
  assign \wptr.add_i  = enq_i;
  assign \wptr.clk  = clk_i;
  assign \wptr.o  = \wptr.ptr_r ;
  assign \wptr.reset_i  = reset_i;
  assign wptr_r = \wptr.ptr_r ;
  assign wptr_r_o = \wptr.ptr_r ;
endmodule
