module bsg_adder_cin(a_i, b_i, cin_i, o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  input [15:0] a_i;
  wire [15:0] a_i;
  input [15:0] b_i;
  wire [15:0] b_i;
  input cin_i;
  wire cin_i;
  output [15:0] o;
  wire [15:0] o;
  assign _035_ = ~(a_i[12] ^ b_i[12]);
  assign _036_ = ~(a_i[11] & b_i[11]);
  assign _037_ = ~(a_i[11] ^ b_i[11]);
  assign _038_ = ~(a_i[10] & b_i[10]);
  assign _039_ = ~(_038_ | _037_);
  assign _040_ = _036_ & ~(_039_);
  assign _041_ = ~(a_i[10] ^ b_i[10]);
  assign _042_ = ~(_041_ | _037_);
  assign _043_ = ~(a_i[9] & b_i[9]);
  assign _044_ = ~(a_i[9] ^ b_i[9]);
  assign _045_ = ~(a_i[8] & b_i[8]);
  assign _046_ = ~(_045_ | _044_);
  assign _047_ = _043_ & ~(_046_);
  assign _048_ = _042_ & ~(_047_);
  assign _049_ = _040_ & ~(_048_);
  assign _050_ = ~(a_i[8] ^ b_i[8]);
  assign _051_ = ~(_050_ | _044_);
  assign _052_ = _051_ & _042_;
  assign _053_ = ~(a_i[7] & b_i[7]);
  assign _054_ = a_i[7] ^ b_i[7];
  assign _055_ = ~(a_i[6] & b_i[6]);
  assign _056_ = _054_ & ~(_055_);
  assign _057_ = _053_ & ~(_056_);
  assign _058_ = ~(a_i[6] ^ b_i[6]);
  assign _059_ = _054_ & ~(_058_);
  assign _060_ = ~(a_i[5] & b_i[5]);
  assign _061_ = ~(a_i[5] ^ b_i[5]);
  assign _062_ = ~(a_i[4] & b_i[4]);
  assign _063_ = ~(_062_ | _061_);
  assign _064_ = _060_ & ~(_063_);
  assign _065_ = _059_ & ~(_064_);
  assign _066_ = _057_ & ~(_065_);
  assign _067_ = ~(a_i[4] ^ b_i[4]);
  assign _068_ = _067_ | _061_;
  assign _069_ = _059_ & ~(_068_);
  assign _070_ = ~(a_i[3] & b_i[3]);
  assign _071_ = a_i[3] ^ b_i[3];
  assign _072_ = ~(a_i[2] & b_i[2]);
  assign _073_ = _071_ & ~(_072_);
  assign _074_ = _070_ & ~(_073_);
  assign _075_ = ~(a_i[2] ^ b_i[2]);
  assign _076_ = _071_ & ~(_075_);
  assign _077_ = ~(a_i[1] & b_i[1]);
  assign _078_ = a_i[1] ^ b_i[1];
  assign _079_ = ~(a_i[0] & b_i[0]);
  assign _080_ = ~(a_i[0] ^ b_i[0]);
  assign _081_ = cin_i & ~(_080_);
  assign _082_ = _079_ & ~(_081_);
  assign _083_ = _078_ & ~(_082_);
  assign _084_ = _077_ & ~(_083_);
  assign _000_ = _076_ & ~(_084_);
  assign _001_ = _074_ & ~(_000_);
  assign _002_ = _069_ & ~(_001_);
  assign _003_ = _066_ & ~(_002_);
  assign _004_ = _052_ & ~(_003_);
  assign _005_ = _049_ & ~(_004_);
  assign o[12] = _005_ ^ _035_;
  assign _006_ = ~(a_i[13] ^ b_i[13]);
  assign _007_ = ~(a_i[12] & b_i[12]);
  assign _008_ = ~(_005_ | _035_);
  assign _009_ = _007_ & ~(_008_);
  assign o[13] = _009_ ^ _006_;
  assign _010_ = ~(a_i[14] ^ b_i[14]);
  assign _011_ = ~(a_i[13] & b_i[13]);
  assign _012_ = ~(_007_ | _006_);
  assign _013_ = _011_ & ~(_012_);
  assign _014_ = _006_ | _035_;
  assign _015_ = ~(_014_ | _005_);
  assign _016_ = _013_ & ~(_015_);
  assign o[14] = _016_ ^ _010_;
  assign _017_ = ~(a_i[15] ^ b_i[15]);
  assign _018_ = ~(a_i[14] & b_i[14]);
  assign _019_ = ~(_016_ | _010_);
  assign _020_ = _018_ & ~(_019_);
  assign o[15] = _020_ ^ _017_;
  assign o[0] = ~(_080_ ^ cin_i);
  assign o[1] = ~(_082_ ^ _078_);
  assign o[2] = _084_ ^ _075_;
  assign _021_ = ~(_084_ | _075_);
  assign _022_ = _021_ | ~(_072_);
  assign o[3] = _022_ ^ _071_;
  assign o[4] = _001_ ^ _067_;
  assign _023_ = ~(_001_ | _067_);
  assign _024_ = _062_ & ~(_023_);
  assign o[5] = _024_ ^ _061_;
  assign _025_ = ~(_001_ | _068_);
  assign _026_ = _064_ & ~(_025_);
  assign o[6] = _026_ ^ _058_;
  assign _027_ = ~(_026_ | _058_);
  assign _028_ = _027_ | ~(_055_);
  assign o[7] = _028_ ^ _054_;
  assign o[8] = _003_ ^ _050_;
  assign _029_ = ~(_003_ | _050_);
  assign _030_ = _045_ & ~(_029_);
  assign o[9] = _030_ ^ _044_;
  assign _031_ = _051_ & ~(_003_);
  assign _032_ = _047_ & ~(_031_);
  assign o[10] = _032_ ^ _041_;
  assign _033_ = ~(_032_ | _041_);
  assign _034_ = _038_ & ~(_033_);
  assign o[11] = _034_ ^ _037_;
endmodule
