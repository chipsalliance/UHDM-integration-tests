module bsg_sbox(clk_i, reset_i, calibration_done_i, channel_active_i, in_v_i, in_data_i, in_yumi_o, in_v_o, in_data_o, in_yumi_i, out_me_v_i, out_me_data_i, out_me_ready_o, out_me_v_o, out_me_data_o, out_me_ready_i);
  wire [4:0] _000_;
  wire [4:0] _001_;
  wire [7:0] _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire [7:0] bk_dpath_sel;
  wire [7:0] bk_dpath_sel_r;
  wire [7:0] bk_sel;
  wire [7:0] bk_sel_r;
  wire [7:0] \bsg.bk_datapath_o ;
  wire [7:0] \bsg.bk_o ;
  wire [7:0] \bsg.fwd_datapath_o ;
  wire [7:0] \bsg.fwd_o ;
  wire [3:0] \bsg.vec_i ;
  input calibration_done_i;
  wire calibration_done_i;
  input [3:0] channel_active_i;
  wire [3:0] channel_active_i;
  input clk_i;
  wire clk_i;
  wire [7:0] fwd_dpath_sel;
  wire [6:0] fwd_dpath_sel_r;
  wire [7:0] fwd_sel;
  reg [7:0] fwd_sel_r;
  input [63:0] in_data_i;
  wire [63:0] in_data_i;
  output [63:0] in_data_o;
  wire [63:0] in_data_o;
  wire [15:0] \in_data_o_int[0] ;
  wire [15:0] \in_data_o_int[1] ;
  wire [15:0] \in_data_o_int[2] ;
  wire [15:0] \in_data_o_int[3] ;
  input [3:0] in_v_i;
  wire [3:0] in_v_i;
  output [3:0] in_v_o;
  wire [3:0] in_v_o;
  wire [3:0] in_v_o_int;
  input [3:0] in_yumi_i;
  wire [3:0] in_yumi_i;
  wire [3:0] in_yumi_i_int;
  output [3:0] in_yumi_o;
  wire [3:0] in_yumi_o;
  input [63:0] out_me_data_i;
  wire [63:0] out_me_data_i;
  wire [15:0] \out_me_data_i_int[0] ;
  wire [15:0] \out_me_data_i_int[1] ;
  wire [15:0] \out_me_data_i_int[2] ;
  wire [15:0] \out_me_data_i_int[3] ;
  output [63:0] out_me_data_o;
  wire [63:0] out_me_data_o;
  input [3:0] out_me_ready_i;
  wire [3:0] out_me_ready_i;
  output [3:0] out_me_ready_o;
  wire [3:0] out_me_ready_o;
  wire [3:0] out_me_ready_o_int;
  input [3:0] out_me_v_i;
  wire [3:0] out_me_v_i;
  wire [3:0] out_me_v_i_int;
  output [3:0] out_me_v_o;
  wire [3:0] out_me_v_o;
  input reset_i;
  wire reset_i;
  wire [15:0] \sbox[0].backward[0] ;
  reg [3:0] \sbox[0].fi1hot.fwd_sel_one_hot_r ;
  wire [15:0] \sbox[0].forward[0] ;
  wire [15:0] \sbox[0].forward[1] ;
  wire [15:0] \sbox[0].forward[2] ;
  wire [15:0] \sbox[0].forward[3] ;
  wire [15:0] \sbox[1].backward[0] ;
  wire [15:0] \sbox[1].backward[1] ;
  wire [7:0] \sbox[1].fi1hot.fwd_sel_one_hot_r ;
  wire [15:0] \sbox[1].forward[0] ;
  wire [15:0] \sbox[1].forward[1] ;
  wire [15:0] \sbox[1].forward[2] ;
  wire [15:0] \sbox[2].backward[0] ;
  wire [15:0] \sbox[2].backward[1] ;
  wire [15:0] \sbox[2].backward[2] ;
  wire [15:0] \sbox[2].fi1hot.fwd_sel_one_hot_r ;
  wire [15:0] \sbox[2].forward[0] ;
  wire [15:0] \sbox[2].forward[1] ;
  wire [15:0] \sbox[3].backward[0] ;
  wire [15:0] \sbox[3].backward[1] ;
  wire [15:0] \sbox[3].backward[2] ;
  wire [15:0] \sbox[3].backward[3] ;
  wire [15:0] \sbox[3].fi1hot.fwd_sel_one_hot_r ;
  wire [15:0] \sbox[3].forward[0] ;
  assign _007_ = \sbox[0].fi1hot.fwd_sel_one_hot_r [0] & in_v_i[0];
  assign _008_ = \sbox[0].fi1hot.fwd_sel_one_hot_r [1] & in_v_i[1];
  assign _009_ = _008_ | _007_;
  assign _010_ = \sbox[0].fi1hot.fwd_sel_one_hot_r [2] & in_v_i[2];
  assign _011_ = \sbox[0].fi1hot.fwd_sel_one_hot_r [3] & in_v_i[3];
  assign _012_ = _011_ | _010_;
  assign in_v_o[0] = _012_ | _009_;
  assign _013_ = \sbox[1].fi1hot.fwd_sel_one_hot_r [4] & in_v_i[0];
  assign _014_ = \sbox[1].fi1hot.fwd_sel_one_hot_r [5] & in_v_i[1];
  assign _015_ = _014_ | _013_;
  assign _016_ = \sbox[1].fi1hot.fwd_sel_one_hot_r [6] & in_v_i[2];
  assign _017_ = \sbox[1].fi1hot.fwd_sel_one_hot_r [7] & in_v_i[3];
  assign _018_ = _017_ | _016_;
  assign in_v_o[1] = _018_ | _015_;
  assign _019_ = \sbox[2].fi1hot.fwd_sel_one_hot_r [8] & in_v_i[0];
  assign _020_ = \sbox[2].fi1hot.fwd_sel_one_hot_r [9] & in_v_i[1];
  assign _021_ = _020_ | _019_;
  assign _022_ = \sbox[2].fi1hot.fwd_sel_one_hot_r [10] & in_v_i[2];
  assign _023_ = \sbox[2].fi1hot.fwd_sel_one_hot_r [11] & in_v_i[3];
  assign _024_ = _023_ | _022_;
  assign in_v_o[2] = _024_ | _021_;
  assign _025_ = \sbox[3].fi1hot.fwd_sel_one_hot_r [12] & in_v_i[0];
  assign _026_ = \sbox[3].fi1hot.fwd_sel_one_hot_r [13] & in_v_i[1];
  assign _027_ = _026_ | _025_;
  assign _028_ = \sbox[3].fi1hot.fwd_sel_one_hot_r [14] & in_v_i[2];
  assign _029_ = \sbox[3].fi1hot.fwd_sel_one_hot_r [15] & in_v_i[3];
  assign _030_ = _029_ | _028_;
  assign in_v_o[3] = _030_ | _027_;
  assign _031_ = ~(bk_dpath_sel_r[6] | bk_dpath_sel_r[7]);
  assign _032_ = ~(bk_dpath_sel_r[6] & bk_dpath_sel_r[7]);
  assign _033_ = out_me_data_i[48] & ~(_032_);
  assign _034_ = bk_dpath_sel_r[6] | ~(bk_dpath_sel_r[7]);
  assign _035_ = out_me_data_i[32] & ~(_034_);
  assign _036_ = _035_ | _033_;
  assign _037_ = bk_dpath_sel_r[7] | ~(bk_dpath_sel_r[6]);
  assign _038_ = out_me_data_i[16] & ~(_037_);
  assign _039_ = _038_ | _036_;
  assign out_me_data_o[48] = _031_ ? out_me_data_i[0] : _039_;
  assign _040_ = out_me_data_i[49] & ~(_032_);
  assign _041_ = out_me_data_i[33] & ~(_034_);
  assign _042_ = _041_ | _040_;
  assign _043_ = out_me_data_i[17] & ~(_037_);
  assign _044_ = _043_ | _042_;
  assign out_me_data_o[49] = _031_ ? out_me_data_i[1] : _044_;
  assign _045_ = out_me_data_i[50] & ~(_032_);
  assign _046_ = out_me_data_i[34] & ~(_034_);
  assign _047_ = _046_ | _045_;
  assign _048_ = out_me_data_i[18] & ~(_037_);
  assign _049_ = _048_ | _047_;
  assign out_me_data_o[50] = _031_ ? out_me_data_i[2] : _049_;
  assign _050_ = out_me_data_i[51] & ~(_032_);
  assign _051_ = out_me_data_i[35] & ~(_034_);
  assign _052_ = _051_ | _050_;
  assign _053_ = out_me_data_i[19] & ~(_037_);
  assign _054_ = _053_ | _052_;
  assign out_me_data_o[51] = _031_ ? out_me_data_i[3] : _054_;
  assign _055_ = out_me_data_i[52] & ~(_032_);
  assign _056_ = out_me_data_i[36] & ~(_034_);
  assign _057_ = _056_ | _055_;
  assign _058_ = out_me_data_i[20] & ~(_037_);
  assign _059_ = _058_ | _057_;
  assign out_me_data_o[52] = _031_ ? out_me_data_i[4] : _059_;
  assign _060_ = out_me_data_i[53] & ~(_032_);
  assign _061_ = out_me_data_i[37] & ~(_034_);
  assign _062_ = _061_ | _060_;
  assign _063_ = out_me_data_i[21] & ~(_037_);
  assign _064_ = _063_ | _062_;
  assign out_me_data_o[53] = _031_ ? out_me_data_i[5] : _064_;
  assign _065_ = out_me_data_i[54] & ~(_032_);
  assign _066_ = out_me_data_i[38] & ~(_034_);
  assign _067_ = _066_ | _065_;
  assign _068_ = out_me_data_i[22] & ~(_037_);
  assign _069_ = _068_ | _067_;
  assign out_me_data_o[54] = _031_ ? out_me_data_i[6] : _069_;
  assign _070_ = out_me_data_i[55] & ~(_032_);
  assign _071_ = out_me_data_i[39] & ~(_034_);
  assign _072_ = _071_ | _070_;
  assign _073_ = out_me_data_i[23] & ~(_037_);
  assign _074_ = _073_ | _072_;
  assign out_me_data_o[55] = _031_ ? out_me_data_i[7] : _074_;
  assign _075_ = out_me_data_i[56] & ~(_032_);
  assign _076_ = out_me_data_i[40] & ~(_034_);
  assign _077_ = _076_ | _075_;
  assign _078_ = out_me_data_i[24] & ~(_037_);
  assign _079_ = _078_ | _077_;
  assign out_me_data_o[56] = _031_ ? out_me_data_i[8] : _079_;
  assign _080_ = out_me_data_i[57] & ~(_032_);
  assign _081_ = out_me_data_i[41] & ~(_034_);
  assign _082_ = _081_ | _080_;
  assign _083_ = out_me_data_i[25] & ~(_037_);
  assign _084_ = _083_ | _082_;
  assign out_me_data_o[57] = _031_ ? out_me_data_i[9] : _084_;
  assign _085_ = out_me_data_i[58] & ~(_032_);
  assign _086_ = out_me_data_i[42] & ~(_034_);
  assign _087_ = _086_ | _085_;
  assign _088_ = out_me_data_i[26] & ~(_037_);
  assign _089_ = _088_ | _087_;
  assign out_me_data_o[58] = _031_ ? out_me_data_i[10] : _089_;
  assign _090_ = out_me_data_i[59] & ~(_032_);
  assign _091_ = out_me_data_i[43] & ~(_034_);
  assign _092_ = _091_ | _090_;
  assign _093_ = out_me_data_i[27] & ~(_037_);
  assign _094_ = _093_ | _092_;
  assign out_me_data_o[59] = _031_ ? out_me_data_i[11] : _094_;
  assign _095_ = out_me_data_i[60] & ~(_032_);
  assign _096_ = out_me_data_i[44] & ~(_034_);
  assign _097_ = _096_ | _095_;
  assign _098_ = out_me_data_i[28] & ~(_037_);
  assign _099_ = _098_ | _097_;
  assign out_me_data_o[60] = _031_ ? out_me_data_i[12] : _099_;
  assign _100_ = out_me_data_i[61] & ~(_032_);
  assign _101_ = out_me_data_i[45] & ~(_034_);
  assign _102_ = _101_ | _100_;
  assign _103_ = out_me_data_i[29] & ~(_037_);
  assign _104_ = _103_ | _102_;
  assign out_me_data_o[61] = _031_ ? out_me_data_i[13] : _104_;
  assign _105_ = out_me_data_i[62] & ~(_032_);
  assign _106_ = out_me_data_i[46] & ~(_034_);
  assign _107_ = _106_ | _105_;
  assign _108_ = out_me_data_i[30] & ~(_037_);
  assign _109_ = _108_ | _107_;
  assign out_me_data_o[62] = _031_ ? out_me_data_i[14] : _109_;
  assign _110_ = out_me_data_i[63] & ~(_032_);
  assign _111_ = out_me_data_i[47] & ~(_034_);
  assign _112_ = _111_ | _110_;
  assign _113_ = out_me_data_i[31] & ~(_037_);
  assign _114_ = _113_ | _112_;
  assign out_me_data_o[63] = _031_ ? out_me_data_i[15] : _114_;
  assign _115_ = bk_dpath_sel_r[4] | ~(bk_dpath_sel_r[5]);
  assign _116_ = bk_dpath_sel_r[5] | ~(bk_dpath_sel_r[4]);
  assign _117_ = _116_ & _115_;
  assign _118_ = out_me_data_i[32] & ~(_115_);
  assign _119_ = out_me_data_i[16] & ~(_116_);
  assign _120_ = _119_ | _118_;
  assign out_me_data_o[32] = _117_ ? out_me_data_i[0] : _120_;
  assign _121_ = out_me_data_i[33] & ~(_115_);
  assign _122_ = out_me_data_i[17] & ~(_116_);
  assign _123_ = _122_ | _121_;
  assign out_me_data_o[33] = _117_ ? out_me_data_i[1] : _123_;
  assign _124_ = out_me_data_i[34] & ~(_115_);
  assign _125_ = out_me_data_i[18] & ~(_116_);
  assign _126_ = _125_ | _124_;
  assign out_me_data_o[34] = _117_ ? out_me_data_i[2] : _126_;
  assign _127_ = out_me_data_i[35] & ~(_115_);
  assign _128_ = out_me_data_i[19] & ~(_116_);
  assign _129_ = _128_ | _127_;
  assign out_me_data_o[35] = _117_ ? out_me_data_i[3] : _129_;
  assign _130_ = out_me_data_i[36] & ~(_115_);
  assign _131_ = out_me_data_i[20] & ~(_116_);
  assign _132_ = _131_ | _130_;
  assign out_me_data_o[36] = _117_ ? out_me_data_i[4] : _132_;
  assign _133_ = out_me_data_i[37] & ~(_115_);
  assign _134_ = out_me_data_i[21] & ~(_116_);
  assign _135_ = _134_ | _133_;
  assign out_me_data_o[37] = _117_ ? out_me_data_i[5] : _135_;
  assign _136_ = out_me_data_i[38] & ~(_115_);
  assign _137_ = out_me_data_i[22] & ~(_116_);
  assign _138_ = _137_ | _136_;
  assign out_me_data_o[38] = _117_ ? out_me_data_i[6] : _138_;
  assign _139_ = out_me_data_i[39] & ~(_115_);
  assign _140_ = out_me_data_i[23] & ~(_116_);
  assign _141_ = _140_ | _139_;
  assign out_me_data_o[39] = _117_ ? out_me_data_i[7] : _141_;
  assign _142_ = out_me_data_i[40] & ~(_115_);
  assign _143_ = out_me_data_i[24] & ~(_116_);
  assign _144_ = _143_ | _142_;
  assign out_me_data_o[40] = _117_ ? out_me_data_i[8] : _144_;
  assign _145_ = out_me_data_i[41] & ~(_115_);
  assign _146_ = out_me_data_i[25] & ~(_116_);
  assign _147_ = _146_ | _145_;
  assign out_me_data_o[41] = _117_ ? out_me_data_i[9] : _147_;
  assign _148_ = out_me_data_i[42] & ~(_115_);
  assign _149_ = out_me_data_i[26] & ~(_116_);
  assign _150_ = _149_ | _148_;
  assign out_me_data_o[42] = _117_ ? out_me_data_i[10] : _150_;
  assign _151_ = out_me_data_i[43] & ~(_115_);
  assign _152_ = out_me_data_i[27] & ~(_116_);
  assign _153_ = _152_ | _151_;
  assign out_me_data_o[43] = _117_ ? out_me_data_i[11] : _153_;
  assign _154_ = out_me_data_i[44] & ~(_115_);
  assign _155_ = out_me_data_i[28] & ~(_116_);
  assign _156_ = _155_ | _154_;
  assign out_me_data_o[44] = _117_ ? out_me_data_i[12] : _156_;
  assign _157_ = out_me_data_i[45] & ~(_115_);
  assign _158_ = out_me_data_i[29] & ~(_116_);
  assign _159_ = _158_ | _157_;
  assign out_me_data_o[45] = _117_ ? out_me_data_i[13] : _159_;
  assign _160_ = out_me_data_i[46] & ~(_115_);
  assign _161_ = out_me_data_i[30] & ~(_116_);
  assign _162_ = _161_ | _160_;
  assign out_me_data_o[46] = _117_ ? out_me_data_i[14] : _162_;
  assign _163_ = out_me_data_i[47] & ~(_115_);
  assign _164_ = out_me_data_i[31] & ~(_116_);
  assign _165_ = _164_ | _163_;
  assign out_me_data_o[47] = _117_ ? out_me_data_i[15] : _165_;
  assign _166_ = bk_dpath_sel_r[4] | ~(fwd_dpath_sel_r[3]);
  assign _167_ = fwd_dpath_sel_r[3] | ~(bk_dpath_sel_r[4]);
  assign _168_ = _167_ & _166_;
  assign _169_ = in_data_i[48] & ~(_166_);
  assign _170_ = in_data_i[32] & ~(_167_);
  assign _171_ = _170_ | _169_;
  assign in_data_o[16] = _168_ ? in_data_i[16] : _171_;
  assign _172_ = in_data_i[49] & ~(_166_);
  assign _173_ = in_data_i[33] & ~(_167_);
  assign _174_ = _173_ | _172_;
  assign in_data_o[17] = _168_ ? in_data_i[17] : _174_;
  assign _175_ = in_data_i[50] & ~(_166_);
  assign _176_ = in_data_i[34] & ~(_167_);
  assign _177_ = _176_ | _175_;
  assign in_data_o[18] = _168_ ? in_data_i[18] : _177_;
  assign _178_ = in_data_i[51] & ~(_166_);
  assign _179_ = in_data_i[35] & ~(_167_);
  assign _180_ = _179_ | _178_;
  assign in_data_o[19] = _168_ ? in_data_i[19] : _180_;
  assign _181_ = in_data_i[52] & ~(_166_);
  assign _182_ = in_data_i[36] & ~(_167_);
  assign _183_ = _182_ | _181_;
  assign in_data_o[20] = _168_ ? in_data_i[20] : _183_;
  assign _184_ = in_data_i[53] & ~(_166_);
  assign _185_ = in_data_i[37] & ~(_167_);
  assign _186_ = _185_ | _184_;
  assign in_data_o[21] = _168_ ? in_data_i[21] : _186_;
  assign _187_ = in_data_i[54] & ~(_166_);
  assign _188_ = in_data_i[38] & ~(_167_);
  assign _189_ = _188_ | _187_;
  assign in_data_o[22] = _168_ ? in_data_i[22] : _189_;
  assign _190_ = in_data_i[55] & ~(_166_);
  assign _191_ = in_data_i[39] & ~(_167_);
  assign _192_ = _191_ | _190_;
  assign in_data_o[23] = _168_ ? in_data_i[23] : _192_;
  assign _193_ = in_data_i[56] & ~(_166_);
  assign _194_ = in_data_i[40] & ~(_167_);
  assign _195_ = _194_ | _193_;
  assign in_data_o[24] = _168_ ? in_data_i[24] : _195_;
  assign _196_ = in_data_i[57] & ~(_166_);
  assign _197_ = in_data_i[41] & ~(_167_);
  assign _198_ = _197_ | _196_;
  assign in_data_o[25] = _168_ ? in_data_i[25] : _198_;
  assign _199_ = in_data_i[58] & ~(_166_);
  assign _200_ = in_data_i[42] & ~(_167_);
  assign _201_ = _200_ | _199_;
  assign in_data_o[26] = _168_ ? in_data_i[26] : _201_;
  assign _202_ = in_data_i[59] & ~(_166_);
  assign _203_ = in_data_i[43] & ~(_167_);
  assign _204_ = _203_ | _202_;
  assign in_data_o[27] = _168_ ? in_data_i[27] : _204_;
  assign _205_ = in_data_i[60] & ~(_166_);
  assign _206_ = in_data_i[44] & ~(_167_);
  assign _207_ = _206_ | _205_;
  assign in_data_o[28] = _168_ ? in_data_i[28] : _207_;
  assign _208_ = in_data_i[61] & ~(_166_);
  assign _209_ = in_data_i[45] & ~(_167_);
  assign _210_ = _209_ | _208_;
  assign in_data_o[29] = _168_ ? in_data_i[29] : _210_;
  assign _211_ = in_data_i[62] & ~(_166_);
  assign _212_ = in_data_i[46] & ~(_167_);
  assign _213_ = _212_ | _211_;
  assign in_data_o[30] = _168_ ? in_data_i[30] : _213_;
  assign _214_ = in_data_i[63] & ~(_166_);
  assign _215_ = in_data_i[47] & ~(_167_);
  assign _216_ = _215_ | _214_;
  assign in_data_o[31] = _168_ ? in_data_i[31] : _216_;
  assign _217_ = ~(fwd_dpath_sel_r[0] | fwd_dpath_sel_r[1]);
  assign _218_ = ~(fwd_dpath_sel_r[0] & fwd_dpath_sel_r[1]);
  assign _219_ = in_data_i[48] & ~(_218_);
  assign _220_ = fwd_dpath_sel_r[0] | ~(fwd_dpath_sel_r[1]);
  assign _221_ = in_data_i[32] & ~(_220_);
  assign _222_ = _221_ | _219_;
  assign _223_ = fwd_dpath_sel_r[1] | ~(fwd_dpath_sel_r[0]);
  assign _224_ = in_data_i[16] & ~(_223_);
  assign _225_ = _224_ | _222_;
  assign in_data_o[0] = _217_ ? in_data_i[0] : _225_;
  assign _226_ = in_data_i[49] & ~(_218_);
  assign _227_ = in_data_i[33] & ~(_220_);
  assign _228_ = _227_ | _226_;
  assign _229_ = in_data_i[17] & ~(_223_);
  assign _230_ = _229_ | _228_;
  assign in_data_o[1] = _217_ ? in_data_i[1] : _230_;
  assign _231_ = in_data_i[50] & ~(_218_);
  assign _232_ = in_data_i[34] & ~(_220_);
  assign _233_ = _232_ | _231_;
  assign _234_ = in_data_i[18] & ~(_223_);
  assign _235_ = _234_ | _233_;
  assign in_data_o[2] = _217_ ? in_data_i[2] : _235_;
  assign _236_ = in_data_i[51] & ~(_218_);
  assign _237_ = in_data_i[35] & ~(_220_);
  assign _238_ = _237_ | _236_;
  assign _239_ = in_data_i[19] & ~(_223_);
  assign _240_ = _239_ | _238_;
  assign in_data_o[3] = _217_ ? in_data_i[3] : _240_;
  assign _241_ = in_data_i[52] & ~(_218_);
  assign _242_ = in_data_i[36] & ~(_220_);
  assign _243_ = _242_ | _241_;
  assign _244_ = in_data_i[20] & ~(_223_);
  assign _245_ = _244_ | _243_;
  assign in_data_o[4] = _217_ ? in_data_i[4] : _245_;
  assign _246_ = in_data_i[53] & ~(_218_);
  assign _247_ = in_data_i[37] & ~(_220_);
  assign _248_ = _247_ | _246_;
  assign _249_ = in_data_i[21] & ~(_223_);
  assign _250_ = _249_ | _248_;
  assign in_data_o[5] = _217_ ? in_data_i[5] : _250_;
  assign _251_ = in_data_i[54] & ~(_218_);
  assign _252_ = in_data_i[38] & ~(_220_);
  assign _253_ = _252_ | _251_;
  assign _254_ = in_data_i[22] & ~(_223_);
  assign _255_ = _254_ | _253_;
  assign in_data_o[6] = _217_ ? in_data_i[6] : _255_;
  assign _256_ = in_data_i[55] & ~(_218_);
  assign _257_ = in_data_i[39] & ~(_220_);
  assign _258_ = _257_ | _256_;
  assign _259_ = in_data_i[23] & ~(_223_);
  assign _260_ = _259_ | _258_;
  assign in_data_o[7] = _217_ ? in_data_i[7] : _260_;
  assign _261_ = in_data_i[56] & ~(_218_);
  assign _262_ = in_data_i[40] & ~(_220_);
  assign _263_ = _262_ | _261_;
  assign _264_ = in_data_i[24] & ~(_223_);
  assign _265_ = _264_ | _263_;
  assign in_data_o[8] = _217_ ? in_data_i[8] : _265_;
  assign _266_ = in_data_i[57] & ~(_218_);
  assign _267_ = in_data_i[41] & ~(_220_);
  assign _268_ = _267_ | _266_;
  assign _269_ = in_data_i[25] & ~(_223_);
  assign _270_ = _269_ | _268_;
  assign in_data_o[9] = _217_ ? in_data_i[9] : _270_;
  assign _271_ = in_data_i[58] & ~(_218_);
  assign _272_ = in_data_i[42] & ~(_220_);
  assign _273_ = _272_ | _271_;
  assign _274_ = in_data_i[26] & ~(_223_);
  assign _275_ = _274_ | _273_;
  assign in_data_o[10] = _217_ ? in_data_i[10] : _275_;
  assign _276_ = in_data_i[59] & ~(_218_);
  assign _277_ = in_data_i[43] & ~(_220_);
  assign _278_ = _277_ | _276_;
  assign _279_ = in_data_i[27] & ~(_223_);
  assign _280_ = _279_ | _278_;
  assign in_data_o[11] = _217_ ? in_data_i[11] : _280_;
  assign _281_ = in_data_i[60] & ~(_218_);
  assign _282_ = in_data_i[44] & ~(_220_);
  assign _283_ = _282_ | _281_;
  assign _284_ = in_data_i[28] & ~(_223_);
  assign _285_ = _284_ | _283_;
  assign in_data_o[12] = _217_ ? in_data_i[12] : _285_;
  assign _286_ = in_data_i[61] & ~(_218_);
  assign _287_ = in_data_i[45] & ~(_220_);
  assign _288_ = _287_ | _286_;
  assign _289_ = in_data_i[29] & ~(_223_);
  assign _290_ = _289_ | _288_;
  assign in_data_o[13] = _217_ ? in_data_i[13] : _290_;
  assign _291_ = in_data_i[62] & ~(_218_);
  assign _292_ = in_data_i[46] & ~(_220_);
  assign _293_ = _292_ | _291_;
  assign _294_ = in_data_i[30] & ~(_223_);
  assign _295_ = _294_ | _293_;
  assign in_data_o[14] = _217_ ? in_data_i[14] : _295_;
  assign _296_ = in_data_i[63] & ~(_218_);
  assign _297_ = in_data_i[47] & ~(_220_);
  assign _298_ = _297_ | _296_;
  assign _299_ = in_data_i[31] & ~(_223_);
  assign _300_ = _299_ | _298_;
  assign in_data_o[15] = _217_ ? in_data_i[15] : _300_;
  assign _002_[1] = ~channel_active_i[0];
  assign _301_ = ~channel_active_i[2];
  assign _002_[2] = channel_active_i[0] | ~(channel_active_i[1]);
  assign _346_ = channel_active_i[2] ? _002_[2] : channel_active_i[0];
  assign fwd_sel[0] = ~_346_;
  assign _302_ = channel_active_i[2] & ~(_002_[2]);
  assign _303_ = _301_ & ~(_002_[2]);
  assign _304_ = _303_ | _302_;
  assign _000_[0] = channel_active_i[3] ? fwd_sel[0] : _304_;
  assign fwd_sel[1] = ~(channel_active_i[1] | channel_active_i[0]);
  assign _305_ = fwd_sel[1] & ~(_301_);
  assign _000_[1] = channel_active_i[3] ? fwd_sel[1] : _305_;
  assign _306_ = ~(channel_active_i[1] & channel_active_i[0]);
  assign _001_[2] = channel_active_i[2] & ~(_306_);
  assign _307_ = channel_active_i[1] & channel_active_i[0];
  assign _308_ = channel_active_i[1] | channel_active_i[0];
  assign _006_ = channel_active_i[2] ? _308_ : _307_;
  assign _309_ = _301_ & ~(_306_);
  assign _310_ = _309_ | _001_[2];
  assign _001_[0] = channel_active_i[3] ? _307_ : _310_;
  assign fwd_sel[3] = ~_307_;
  assign _311_ = channel_active_i[1] ^ channel_active_i[0];
  assign _000_[2] = _311_ & ~(_301_);
  assign _003_ = channel_active_i[2] ? fwd_sel[1] : _311_;
  assign _004_ = channel_active_i[2] ? _311_ : _307_;
  assign _002_[5] = _307_ | _301_;
  assign _312_ = _307_ | fwd_sel[1];
  assign _005_ = channel_active_i[2] ? _312_ : _311_;
  assign _002_[4] = _311_ | _301_;
  assign _002_[3] = ~channel_active_i[1];
  assign out_me_data_o[16] = bk_dpath_sel_r[2] ? out_me_data_i[16] : out_me_data_i[0];
  assign out_me_data_o[17] = bk_dpath_sel_r[2] ? out_me_data_i[17] : out_me_data_i[1];
  assign out_me_data_o[18] = bk_dpath_sel_r[2] ? out_me_data_i[18] : out_me_data_i[2];
  assign out_me_data_o[19] = bk_dpath_sel_r[2] ? out_me_data_i[19] : out_me_data_i[3];
  assign out_me_data_o[20] = bk_dpath_sel_r[2] ? out_me_data_i[20] : out_me_data_i[4];
  assign out_me_data_o[21] = bk_dpath_sel_r[2] ? out_me_data_i[21] : out_me_data_i[5];
  assign out_me_data_o[22] = bk_dpath_sel_r[2] ? out_me_data_i[22] : out_me_data_i[6];
  assign out_me_data_o[23] = bk_dpath_sel_r[2] ? out_me_data_i[23] : out_me_data_i[7];
  assign out_me_data_o[24] = bk_dpath_sel_r[2] ? out_me_data_i[24] : out_me_data_i[8];
  assign out_me_data_o[25] = bk_dpath_sel_r[2] ? out_me_data_i[25] : out_me_data_i[9];
  assign out_me_data_o[26] = bk_dpath_sel_r[2] ? out_me_data_i[26] : out_me_data_i[10];
  assign out_me_data_o[27] = bk_dpath_sel_r[2] ? out_me_data_i[27] : out_me_data_i[11];
  assign out_me_data_o[28] = bk_dpath_sel_r[2] ? out_me_data_i[28] : out_me_data_i[12];
  assign out_me_data_o[29] = bk_dpath_sel_r[2] ? out_me_data_i[29] : out_me_data_i[13];
  assign out_me_data_o[30] = bk_dpath_sel_r[2] ? out_me_data_i[30] : out_me_data_i[14];
  assign out_me_data_o[31] = bk_dpath_sel_r[2] ? out_me_data_i[31] : out_me_data_i[15];
  assign _313_ = ~channel_active_i[3];
  assign _314_ = _312_ | _301_;
  assign _315_ = channel_active_i[2] ? _312_ : _308_;
  assign fwd_sel[2] = channel_active_i[3] ? _315_ : _314_;
  assign _316_ = _307_ & ~(_301_);
  assign _317_ = channel_active_i[2] ? _307_ : _306_;
  assign _348_ = channel_active_i[3] ? _317_ : _316_;
  assign fwd_sel[4] = ~_348_;
  assign _318_ = _308_ | _301_;
  assign fwd_sel[5] = _318_ | _313_;
  assign _319_ = _002_[2] & ~(_301_);
  assign _349_ = channel_active_i[3] & ~(_319_);
  assign fwd_sel[6] = ~_349_;
  assign fwd_sel[7] = _002_[5] | _313_;
  assign in_data_o[32] = fwd_dpath_sel_r[4] ? in_data_i[48] : in_data_i[32];
  assign in_data_o[33] = fwd_dpath_sel_r[4] ? in_data_i[49] : in_data_i[33];
  assign in_data_o[34] = fwd_dpath_sel_r[4] ? in_data_i[50] : in_data_i[34];
  assign in_data_o[35] = fwd_dpath_sel_r[4] ? in_data_i[51] : in_data_i[35];
  assign in_data_o[36] = fwd_dpath_sel_r[4] ? in_data_i[52] : in_data_i[36];
  assign in_data_o[37] = fwd_dpath_sel_r[4] ? in_data_i[53] : in_data_i[37];
  assign in_data_o[38] = fwd_dpath_sel_r[4] ? in_data_i[54] : in_data_i[38];
  assign in_data_o[39] = fwd_dpath_sel_r[4] ? in_data_i[55] : in_data_i[39];
  assign in_data_o[40] = fwd_dpath_sel_r[4] ? in_data_i[56] : in_data_i[40];
  assign in_data_o[41] = fwd_dpath_sel_r[4] ? in_data_i[57] : in_data_i[41];
  assign in_data_o[42] = fwd_dpath_sel_r[4] ? in_data_i[58] : in_data_i[42];
  assign in_data_o[43] = fwd_dpath_sel_r[4] ? in_data_i[59] : in_data_i[43];
  assign in_data_o[44] = fwd_dpath_sel_r[4] ? in_data_i[60] : in_data_i[44];
  assign in_data_o[45] = fwd_dpath_sel_r[4] ? in_data_i[61] : in_data_i[45];
  assign in_data_o[46] = fwd_dpath_sel_r[4] ? in_data_i[62] : in_data_i[46];
  assign in_data_o[47] = fwd_dpath_sel_r[4] ? in_data_i[63] : in_data_i[47];
  assign _320_ = bk_sel_r[1] ? in_yumi_i[1] : in_yumi_i[0];
  assign _321_ = bk_sel_r[1] ? in_yumi_i[3] : in_yumi_i[2];
  assign in_yumi_o[0] = bk_sel_r[1] ? _321_ : _320_;
  assign _322_ = bk_sel_r[1] ? out_me_v_i[1] : out_me_v_i[0];
  assign _323_ = bk_sel_r[1] ? out_me_v_i[3] : out_me_v_i[2];
  assign out_me_v_o[0] = bk_sel_r[1] ? _323_ : _322_;
  assign _324_ = fwd_sel_r[0] ? out_me_ready_i[1] : out_me_ready_i[0];
  assign _325_ = fwd_sel_r[0] ? out_me_ready_i[3] : out_me_ready_i[2];
  assign out_me_ready_o[0] = fwd_sel_r[1] ? _325_ : _324_;
  assign _326_ = bk_sel_r[2] ? in_yumi_i[1] : in_yumi_i[0];
  assign _327_ = bk_sel_r[2] ? in_yumi_i[3] : in_yumi_i[2];
  assign in_yumi_o[1] = bk_sel_r[3] ? _327_ : _326_;
  assign _328_ = bk_sel_r[2] ? out_me_v_i[1] : out_me_v_i[0];
  assign _329_ = bk_sel_r[2] ? out_me_v_i[3] : out_me_v_i[2];
  assign out_me_v_o[1] = bk_sel_r[3] ? _329_ : _328_;
  assign _330_ = fwd_sel_r[2] ? out_me_ready_i[1] : out_me_ready_i[0];
  assign _331_ = fwd_sel_r[2] ? out_me_ready_i[3] : out_me_ready_i[2];
  assign out_me_ready_o[1] = fwd_sel_r[3] ? _331_ : _330_;
  assign _332_ = bk_sel_r[4] ? in_yumi_i[1] : in_yumi_i[0];
  assign _333_ = bk_sel_r[4] ? in_yumi_i[3] : in_yumi_i[2];
  assign in_yumi_o[2] = bk_sel_r[5] ? _333_ : _332_;
  assign _334_ = bk_sel_r[4] ? out_me_v_i[1] : out_me_v_i[0];
  assign _335_ = bk_sel_r[4] ? out_me_v_i[3] : out_me_v_i[2];
  assign out_me_v_o[2] = bk_sel_r[5] ? _335_ : _334_;
  assign _336_ = fwd_sel_r[4] ? out_me_ready_i[1] : out_me_ready_i[0];
  assign _337_ = fwd_sel_r[4] ? out_me_ready_i[3] : out_me_ready_i[2];
  assign out_me_ready_o[2] = fwd_sel_r[5] ? _337_ : _336_;
  assign _338_ = bk_sel_r[6] ? in_yumi_i[1] : in_yumi_i[0];
  assign _339_ = bk_sel_r[6] ? in_yumi_i[3] : in_yumi_i[2];
  assign in_yumi_o[3] = bk_sel_r[7] ? _339_ : _338_;
  assign _340_ = bk_sel_r[6] ? out_me_v_i[1] : out_me_v_i[0];
  assign _341_ = bk_sel_r[6] ? out_me_v_i[3] : out_me_v_i[2];
  assign out_me_v_o[3] = bk_sel_r[7] ? _341_ : _340_;
  assign _342_ = fwd_sel_r[6] ? out_me_ready_i[1] : out_me_ready_i[0];
  assign _343_ = fwd_sel_r[6] ? out_me_ready_i[3] : out_me_ready_i[2];
  assign out_me_ready_o[3] = fwd_sel_r[7] ? _343_ : _342_;
  assign _344_ = ~(_314_ & _313_);
  assign _345_ = _315_ & ~(_313_);
  assign _347_ = _344_ & ~(_345_);
  always @(posedge clk_i)
    if (!fwd_sel[1]) \sbox[0].fi1hot.fwd_sel_one_hot_r [3] <= 1'h0;
    else \sbox[0].fi1hot.fwd_sel_one_hot_r [3] <= fwd_sel[0];
  reg \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[7] ;
  always @(posedge clk_i)
    if (_307_) \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[7]  <= 1'h0;
    else \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[7]  <= fwd_sel[2];
  assign \sbox[1].fi1hot.fwd_sel_one_hot_r [7] = \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[7] ;
  reg \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[11] ;
  always @(posedge clk_i)
    if (!fwd_sel[5]) \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[11]  <= 1'h0;
    else \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[11]  <= fwd_sel[4];
  assign \sbox[2].fi1hot.fwd_sel_one_hot_r [11] = \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[11] ;
  reg \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[15] ;
  always @(posedge clk_i)
    if (!fwd_sel[7]) \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[15]  <= 1'h0;
    else \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[15]  <= fwd_sel[6];
  assign \sbox[3].fi1hot.fwd_sel_one_hot_r [15] = \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[15] ;
  reg \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[12] ;
  always @(posedge clk_i)
    if (fwd_sel[7]) \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[12]  <= 1'h0;
    else \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[12]  <= _349_;
  assign \sbox[3].fi1hot.fwd_sel_one_hot_r [12] = \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[12] ;
  reg \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[13] ;
  always @(posedge clk_i)
    if (fwd_sel[7]) \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[13]  <= 1'h0;
    else \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[13]  <= fwd_sel[6];
  assign \sbox[3].fi1hot.fwd_sel_one_hot_r [13] = \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[13] ;
  reg \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[14] ;
  always @(posedge clk_i)
    if (!fwd_sel[7]) \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[14]  <= 1'h0;
    else \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[14]  <= _349_;
  assign \sbox[3].fi1hot.fwd_sel_one_hot_r [14] = \sbox_reg[3].fi1hot.fwd_sel_one_hot_r[14] ;
  reg \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[8] ;
  always @(posedge clk_i)
    if (fwd_sel[5]) \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[8]  <= 1'h0;
    else \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[8]  <= _348_;
  assign \sbox[2].fi1hot.fwd_sel_one_hot_r [8] = \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[8] ;
  reg \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[9] ;
  always @(posedge clk_i)
    if (fwd_sel[5]) \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[9]  <= 1'h0;
    else \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[9]  <= fwd_sel[4];
  assign \sbox[2].fi1hot.fwd_sel_one_hot_r [9] = \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[9] ;
  reg \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[10] ;
  always @(posedge clk_i)
    if (!fwd_sel[5]) \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[10]  <= 1'h0;
    else \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[10]  <= _348_;
  assign \sbox[2].fi1hot.fwd_sel_one_hot_r [10] = \sbox_reg[2].fi1hot.fwd_sel_one_hot_r[10] ;
  reg \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[4] ;
  always @(posedge clk_i)
    if (!_307_) \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[4]  <= 1'h0;
    else \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[4]  <= _347_;
  assign \sbox[1].fi1hot.fwd_sel_one_hot_r [4] = \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[4] ;
  reg \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[5] ;
  always @(posedge clk_i)
    if (!_307_) \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[5]  <= 1'h0;
    else \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[5]  <= fwd_sel[2];
  assign \sbox[1].fi1hot.fwd_sel_one_hot_r [5] = \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[5] ;
  reg \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[6] ;
  always @(posedge clk_i)
    if (_307_) \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[6]  <= 1'h0;
    else \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[6]  <= _347_;
  assign \sbox[1].fi1hot.fwd_sel_one_hot_r [6] = \sbox_reg[1].fi1hot.fwd_sel_one_hot_r[6] ;
  always @(posedge clk_i)
    if (fwd_sel[1]) \sbox[0].fi1hot.fwd_sel_one_hot_r [0] <= 1'h0;
    else \sbox[0].fi1hot.fwd_sel_one_hot_r [0] <= _346_;
  always @(posedge clk_i)
    if (fwd_sel[1]) \sbox[0].fi1hot.fwd_sel_one_hot_r [1] <= 1'h0;
    else \sbox[0].fi1hot.fwd_sel_one_hot_r [1] <= fwd_sel[0];
  always @(posedge clk_i)
    if (!fwd_sel[1]) \sbox[0].fi1hot.fwd_sel_one_hot_r [2] <= 1'h0;
    else \sbox[0].fi1hot.fwd_sel_one_hot_r [2] <= _346_;
  reg \fwd_dpath_sel_r_reg[3] ;
  always @(posedge clk_i)
    if (!channel_active_i[3]) \fwd_dpath_sel_r_reg[3]  <= 1'h0;
    else \fwd_dpath_sel_r_reg[3]  <= _003_;
  assign fwd_dpath_sel_r[3] = \fwd_dpath_sel_r_reg[3] ;
  reg \fwd_dpath_sel_r_reg[4] ;
  always @(posedge clk_i)
    if (!channel_active_i[3]) \fwd_dpath_sel_r_reg[4]  <= 1'h0;
    else \fwd_dpath_sel_r_reg[4]  <= _004_;
  assign fwd_dpath_sel_r[4] = \fwd_dpath_sel_r_reg[4] ;
  reg \bk_sel_r_reg[1] ;
  always @(posedge clk_i)
    \bk_sel_r_reg[1]  <= _002_[1];
  assign bk_sel_r[1] = \bk_sel_r_reg[1] ;
  reg \bk_sel_r_reg[2] ;
  always @(posedge clk_i)
    \bk_sel_r_reg[2]  <= _002_[2];
  assign bk_sel_r[2] = \bk_sel_r_reg[2] ;
  reg \bk_sel_r_reg[3] ;
  always @(posedge clk_i)
    \bk_sel_r_reg[3]  <= _002_[3];
  assign bk_sel_r[3] = \bk_sel_r_reg[3] ;
  reg \bk_sel_r_reg[4] ;
  always @(posedge clk_i)
    \bk_sel_r_reg[4]  <= _002_[4];
  assign bk_sel_r[4] = \bk_sel_r_reg[4] ;
  reg \bk_sel_r_reg[5] ;
  always @(posedge clk_i)
    \bk_sel_r_reg[5]  <= _002_[5];
  assign bk_sel_r[5] = \bk_sel_r_reg[5] ;
  reg \bk_sel_r_reg[6] ;
  always @(posedge clk_i)
    if (!channel_active_i[3]) \bk_sel_r_reg[6]  <= 1'h1;
    else \bk_sel_r_reg[6]  <= _005_;
  assign bk_sel_r[6] = \bk_sel_r_reg[6] ;
  reg \bk_sel_r_reg[7] ;
  always @(posedge clk_i)
    if (!channel_active_i[3]) \bk_sel_r_reg[7]  <= 1'h1;
    else \bk_sel_r_reg[7]  <= _006_;
  assign bk_sel_r[7] = \bk_sel_r_reg[7] ;
  always @(posedge clk_i)
    fwd_sel_r[0] <= fwd_sel[0];
  always @(posedge clk_i)
    fwd_sel_r[1] <= fwd_sel[1];
  always @(posedge clk_i)
    fwd_sel_r[2] <= fwd_sel[2];
  always @(posedge clk_i)
    fwd_sel_r[3] <= fwd_sel[3];
  always @(posedge clk_i)
    fwd_sel_r[4] <= fwd_sel[4];
  always @(posedge clk_i)
    fwd_sel_r[5] <= fwd_sel[5];
  always @(posedge clk_i)
    fwd_sel_r[6] <= fwd_sel[6];
  always @(posedge clk_i)
    fwd_sel_r[7] <= fwd_sel[7];
  reg \bk_dpath_sel_r_reg[6] ;
  always @(posedge clk_i)
    if (!channel_active_i[3]) \bk_dpath_sel_r_reg[6]  <= 1'h0;
    else \bk_dpath_sel_r_reg[6]  <= _005_;
  assign bk_dpath_sel_r[6] = \bk_dpath_sel_r_reg[6] ;
  reg \bk_dpath_sel_r_reg[7] ;
  always @(posedge clk_i)
    if (!channel_active_i[3]) \bk_dpath_sel_r_reg[7]  <= 1'h0;
    else \bk_dpath_sel_r_reg[7]  <= _006_;
  assign bk_dpath_sel_r[7] = \bk_dpath_sel_r_reg[7] ;
  reg \bk_dpath_sel_r_reg[2] ;
  always @(posedge clk_i)
    \bk_dpath_sel_r_reg[2]  <= _001_[0];
  assign bk_dpath_sel_r[2] = \bk_dpath_sel_r_reg[2] ;
  reg \bk_dpath_sel_r_reg[4] ;
  always @(posedge clk_i)
    \bk_dpath_sel_r_reg[4]  <= _000_[2];
  assign bk_dpath_sel_r[4] = \bk_dpath_sel_r_reg[4] ;
  reg \bk_dpath_sel_r_reg[5] ;
  always @(posedge clk_i)
    \bk_dpath_sel_r_reg[5]  <= _001_[2];
  assign bk_dpath_sel_r[5] = \bk_dpath_sel_r_reg[5] ;
  reg \fwd_dpath_sel_r_reg[0] ;
  always @(posedge clk_i)
    \fwd_dpath_sel_r_reg[0]  <= _000_[0];
  assign fwd_dpath_sel_r[0] = \fwd_dpath_sel_r_reg[0] ;
  reg \fwd_dpath_sel_r_reg[1] ;
  always @(posedge clk_i)
    \fwd_dpath_sel_r_reg[1]  <= _000_[1];
  assign fwd_dpath_sel_r[1] = \fwd_dpath_sel_r_reg[1] ;
  assign _001_[1] = _000_[2];
  assign _002_[0] = _002_[1];
  assign bk_dpath_sel = 8'bxxxx0x00;
  assign { bk_dpath_sel_r[3], bk_dpath_sel_r[1:0] } = 3'h0;
  assign bk_sel = 8'hxx;
  assign bk_sel_r[0] = bk_sel_r[1];
  assign \bsg.bk_datapath_o  = 8'bxxxx0x00;
  assign \bsg.bk_o  = 8'hxx;
  assign \bsg.fwd_datapath_o  = 8'b000xxxxx;
  assign \bsg.fwd_o  = fwd_sel;
  assign \bsg.vec_i  = channel_active_i;
  assign fwd_dpath_sel = 8'b000xxxxx;
  assign { fwd_dpath_sel_r[6:5], fwd_dpath_sel_r[2] } = { 2'h0, bk_dpath_sel_r[4] };
  assign in_data_o[63:48] = in_data_i[63:48];
  assign \in_data_o_int[0]  = in_data_o[15:0];
  assign \in_data_o_int[1]  = in_data_o[31:16];
  assign \in_data_o_int[2]  = in_data_o[47:32];
  assign \in_data_o_int[3]  = in_data_i[63:48];
  assign in_v_o_int = in_v_o;
  assign in_yumi_i_int = in_yumi_i;
  assign \out_me_data_i_int[0]  = out_me_data_i[15:0];
  assign \out_me_data_i_int[1]  = out_me_data_i[31:16];
  assign \out_me_data_i_int[2]  = out_me_data_i[47:32];
  assign \out_me_data_i_int[3]  = out_me_data_i[63:48];
  assign out_me_data_o[15:0] = out_me_data_i[15:0];
  assign out_me_ready_o_int = out_me_ready_o;
  assign out_me_v_i_int = out_me_v_i;
  assign \sbox[0].backward[0]  = out_me_data_i[15:0];
  assign \sbox[0].forward[0]  = in_data_i[15:0];
  assign \sbox[0].forward[1]  = in_data_i[31:16];
  assign \sbox[0].forward[2]  = in_data_i[47:32];
  assign \sbox[0].forward[3]  = in_data_i[63:48];
  assign \sbox[1].backward[0]  = out_me_data_i[15:0];
  assign \sbox[1].backward[1]  = out_me_data_i[31:16];
  assign \sbox[1].fi1hot.fwd_sel_one_hot_r [3:0] = 4'hx;
  assign \sbox[1].forward[0]  = in_data_i[31:16];
  assign \sbox[1].forward[1]  = in_data_i[47:32];
  assign \sbox[1].forward[2]  = in_data_i[63:48];
  assign \sbox[2].backward[0]  = out_me_data_i[15:0];
  assign \sbox[2].backward[1]  = out_me_data_i[31:16];
  assign \sbox[2].backward[2]  = out_me_data_i[47:32];
  assign { \sbox[2].fi1hot.fwd_sel_one_hot_r [15:12], \sbox[2].fi1hot.fwd_sel_one_hot_r [7:0] } = 12'hxxx;
  assign \sbox[2].forward[0]  = in_data_i[47:32];
  assign \sbox[2].forward[1]  = in_data_i[63:48];
  assign \sbox[3].backward[0]  = out_me_data_i[15:0];
  assign \sbox[3].backward[1]  = out_me_data_i[31:16];
  assign \sbox[3].backward[2]  = out_me_data_i[47:32];
  assign \sbox[3].backward[3]  = out_me_data_i[63:48];
  assign \sbox[3].fi1hot.fwd_sel_one_hot_r [11:0] = 12'hxxx;
  assign \sbox[3].forward[0]  = in_data_i[63:48];
endmodule
