module top;
   parameter int a = '0;
   parameter int b = '1;
   parameter int c = 'x;
   parameter int d = 'z;
endmodule // top
