module bsg_mul_synth(a_i, b_i, o);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  input [15:0] a_i;
  wire [15:0] a_i;
  input [15:0] b_i;
  wire [15:0] b_i;
  output [31:0] o;
  wire [31:0] o;
  assign o[0] = b_i[0] & a_i[0];
  assign _1189_ = a_i[2] & b_i[0];
  assign _1200_ = b_i[1] & a_i[1];
  assign _1210_ = ~(_1200_ ^ _1189_);
  assign _1221_ = b_i[2] & a_i[0];
  assign _1232_ = _1221_ ^ _1210_;
  assign _1243_ = a_i[1] & b_i[0];
  assign _1254_ = b_i[1] & a_i[0];
  assign _1265_ = _1254_ & _1243_;
  assign o[2] = ~(_1265_ ^ _1232_);
  assign _1286_ = a_i[3] & b_i[0];
  assign _1297_ = b_i[1] & a_i[2];
  assign _1307_ = _1297_ ^ _1286_;
  assign _1318_ = b_i[2] & a_i[1];
  assign _1329_ = ~_1318_;
  assign _1340_ = _1329_ ^ _1307_;
  assign _1351_ = ~(_1200_ & _1189_);
  assign _1362_ = _1221_ & ~(_1210_);
  assign _1373_ = _1351_ & ~(_1362_);
  assign _1384_ = ~(_1373_ ^ _1340_);
  assign _1395_ = b_i[3] & a_i[0];
  assign _1406_ = _1395_ ^ _1384_;
  assign _1416_ = _1265_ & ~(_1232_);
  assign o[3] = ~(_1416_ ^ _1406_);
  assign _1437_ = ~(a_i[4] & b_i[0]);
  assign _1448_ = ~(b_i[1] & a_i[3]);
  assign _1459_ = _1448_ ^ _1437_;
  assign _1470_ = ~(b_i[2] & a_i[2]);
  assign _1481_ = _1470_ ^ _1459_;
  assign _1492_ = ~(_1297_ & _1286_);
  assign _1503_ = _1307_ & ~(_1329_);
  assign _1513_ = _1492_ & ~(_1503_);
  assign _1524_ = _1513_ ^ _1481_;
  assign _1535_ = b_i[3] & a_i[1];
  assign _1546_ = b_i[4] & a_i[0];
  assign _0010_ = ~(_1546_ ^ _1535_);
  assign _0021_ = _0010_ ^ _1524_;
  assign _0032_ = ~_0021_;
  assign _0043_ = _1373_ | _1340_;
  assign _0053_ = _1395_ & ~(_1384_);
  assign _0064_ = _0043_ & ~(_0053_);
  assign _0075_ = _0064_ ^ _0032_;
  assign _0086_ = _1416_ & ~(_1406_);
  assign o[4] = ~(_0086_ ^ _0075_);
  assign _0107_ = ~(a_i[5] & b_i[0]);
  assign _0118_ = ~(b_i[1] & a_i[4]);
  assign _0129_ = _0118_ ^ _0107_;
  assign _0139_ = ~(b_i[2] & a_i[3]);
  assign _0150_ = _0139_ ^ _0129_;
  assign _0161_ = _1448_ | _1437_;
  assign _0172_ = _1459_ & ~(_1470_);
  assign _0183_ = _0161_ & ~(_0172_);
  assign _0194_ = _0183_ ^ _0150_;
  assign _0205_ = ~(b_i[3] & a_i[2]);
  assign _0216_ = b_i[4] & a_i[1];
  assign _0226_ = _0216_ ^ _0205_;
  assign _0237_ = b_i[5] & a_i[0];
  assign _0248_ = _0237_ ^ _0226_;
  assign _0259_ = _0248_ ^ _0194_;
  assign _0270_ = _1513_ | _1481_;
  assign _0281_ = _1524_ & ~(_0010_);
  assign _0291_ = _0270_ & ~(_0281_);
  assign _0302_ = _0291_ ^ _0259_;
  assign _0313_ = _1546_ & _1535_;
  assign _0324_ = ~_0313_;
  assign _0335_ = _0324_ ^ _0302_;
  assign _0346_ = _0032_ & ~(_0064_);
  assign _0357_ = _0346_ ^ _0335_;
  assign _0367_ = _0086_ & ~(_0075_);
  assign o[5] = ~(_0367_ ^ _0357_);
  assign _0388_ = ~(a_i[6] & b_i[0]);
  assign _0399_ = ~(b_i[1] & a_i[5]);
  assign _0410_ = _0399_ ^ _0388_;
  assign _0420_ = ~(b_i[2] & a_i[4]);
  assign _0431_ = _0420_ ^ _0410_;
  assign _0442_ = _0118_ | _0107_;
  assign _0453_ = _0129_ & ~(_0139_);
  assign _0464_ = _0442_ & ~(_0453_);
  assign _0475_ = _0464_ ^ _0431_;
  assign _0485_ = ~(b_i[3] & a_i[3]);
  assign _0496_ = b_i[4] & a_i[2];
  assign _0507_ = _0496_ ^ _0485_;
  assign _0518_ = b_i[5] & a_i[1];
  assign _0529_ = _0518_ ^ _0507_;
  assign _0539_ = _0529_ ^ _0475_;
  assign _0550_ = _0183_ | _0150_;
  assign _0561_ = _0194_ & ~(_0248_);
  assign _0572_ = _0550_ & ~(_0561_);
  assign _0582_ = _0572_ ^ _0539_;
  assign _0593_ = _0216_ & ~(_0205_);
  assign _0604_ = _0237_ & ~(_0226_);
  assign _0614_ = ~(_0604_ | _0593_);
  assign _0625_ = b_i[6] & a_i[0];
  assign _0636_ = _0625_ ^ _0614_;
  assign _0646_ = _0636_ ^ _0582_;
  assign _0657_ = ~_0646_;
  assign _0667_ = _0291_ | _0259_;
  assign _0678_ = _0302_ & ~(_0324_);
  assign _0688_ = _0667_ & ~(_0678_);
  assign _0690_ = _0688_ ^ _0657_;
  assign _0691_ = _0346_ & ~(_0335_);
  assign _0692_ = _0691_ ^ _0690_;
  assign _0693_ = _0367_ & ~(_0357_);
  assign o[6] = ~(_0693_ ^ _0692_);
  assign _0694_ = ~(a_i[8] & b_i[0]);
  assign _0695_ = ~(b_i[1] & a_i[7]);
  assign _0696_ = _0695_ ^ _0694_;
  assign _0697_ = ~(b_i[2] & a_i[6]);
  assign _0698_ = _0697_ ^ _0696_;
  assign _0699_ = ~(a_i[7] & b_i[0]);
  assign _0700_ = b_i[1] & a_i[6];
  assign _0701_ = _0699_ | ~(_0700_);
  assign _0702_ = b_i[2] & a_i[5];
  assign _0703_ = _0700_ ^ _0699_;
  assign _0704_ = _0702_ & ~(_0703_);
  assign _0705_ = _0701_ & ~(_0704_);
  assign _0706_ = _0705_ ^ _0698_;
  assign _0707_ = ~(b_i[3] & a_i[5]);
  assign _0708_ = ~(b_i[4] & a_i[4]);
  assign _0709_ = _0708_ ^ _0707_;
  assign _0710_ = ~(b_i[5] & a_i[3]);
  assign _0711_ = _0710_ ^ _0709_;
  assign _0712_ = _0711_ ^ _0706_;
  assign _0713_ = ~(_0703_ ^ _0702_);
  assign _0714_ = _0399_ | _0388_;
  assign _0715_ = _0410_ & ~(_0420_);
  assign _0716_ = _0714_ & ~(_0715_);
  assign _0717_ = _0716_ | ~(_0713_);
  assign _0718_ = b_i[3] & a_i[4];
  assign _0719_ = b_i[4] & a_i[3];
  assign _0720_ = _0719_ ^ _0718_;
  assign _0721_ = b_i[5] & a_i[2];
  assign _0722_ = _0721_ ^ _0720_;
  assign _0723_ = _0716_ ^ _0713_;
  assign _0724_ = _0722_ & ~(_0723_);
  assign _0725_ = _0717_ & ~(_0724_);
  assign _0726_ = _0725_ ^ _0712_;
  assign _0727_ = _0719_ & _0718_;
  assign _0728_ = _0721_ & _0720_;
  assign _0729_ = ~(_0728_ | _0727_);
  assign _0730_ = ~(b_i[6] & a_i[2]);
  assign _0731_ = b_i[7] & a_i[1];
  assign _0732_ = ~(_0731_ ^ _0730_);
  assign _0733_ = b_i[8] & a_i[0];
  assign _0734_ = ~_0733_;
  assign _0735_ = _0734_ ^ _0732_;
  assign _0736_ = _0735_ ^ _0729_;
  assign _0737_ = b_i[6] & a_i[1];
  assign _0738_ = b_i[7] & a_i[0];
  assign _0739_ = _0738_ & _0737_;
  assign _0740_ = ~_0739_;
  assign _0741_ = _0740_ ^ _0736_;
  assign _0742_ = _0741_ ^ _0726_;
  assign _0743_ = ~(_0723_ ^ _0722_);
  assign _0744_ = _0464_ | _0431_;
  assign _0745_ = _0475_ & ~(_0529_);
  assign _0746_ = _0744_ & ~(_0745_);
  assign _0747_ = _0746_ | ~(_0743_);
  assign _0748_ = _0496_ & ~(_0485_);
  assign _0749_ = _0518_ & ~(_0507_);
  assign _0750_ = ~(_0749_ | _0748_);
  assign _0751_ = ~(_0738_ ^ _0737_);
  assign _0752_ = ~(_0751_ ^ _0750_);
  assign _0753_ = _0746_ ^ _0743_;
  assign _0754_ = ~(_0753_ | _0752_);
  assign _0755_ = _0747_ & ~(_0754_);
  assign _0756_ = _0755_ ^ _0742_;
  assign _0757_ = ~(_0751_ | _0750_);
  assign _0758_ = ~_0757_;
  assign _0759_ = _0758_ ^ _0756_;
  assign _0760_ = ~_0759_;
  assign _0761_ = _0753_ ^ _0752_;
  assign _0762_ = _0572_ | _0539_;
  assign _0763_ = _0582_ & ~(_0636_);
  assign _0764_ = _0762_ & ~(_0763_);
  assign _0765_ = _0764_ | ~(_0761_);
  assign _0766_ = _0625_ & ~(_0614_);
  assign _0767_ = _0764_ ^ _0761_;
  assign _0768_ = _0766_ & ~(_0767_);
  assign _0769_ = _0765_ & ~(_0768_);
  assign _0770_ = _0769_ ^ _0760_;
  assign _0771_ = _0767_ ^ _0766_;
  assign _0772_ = _0657_ & ~(_0688_);
  assign _0773_ = _0772_ & ~(_0771_);
  assign _0774_ = _0773_ ^ _0770_;
  assign _0775_ = _0772_ ^ _0771_;
  assign _0776_ = _0690_ | ~(_0691_);
  assign _0777_ = _0776_ | _0775_;
  assign _0778_ = ~(_0777_ ^ _0774_);
  assign _0779_ = ~(_0776_ ^ _0775_);
  assign _0780_ = _0693_ & ~(_0692_);
  assign _0781_ = _0780_ & ~(_0779_);
  assign _0782_ = ~_0781_;
  assign o[8] = _0782_ ^ _0778_;
  assign _0783_ = ~(a_i[9] & b_i[0]);
  assign _0784_ = ~(b_i[1] & a_i[8]);
  assign _0785_ = _0784_ ^ _0783_;
  assign _0786_ = ~(b_i[2] & a_i[7]);
  assign _0787_ = _0786_ ^ _0785_;
  assign _0788_ = _0695_ | _0694_;
  assign _0789_ = _0696_ & ~(_0697_);
  assign _0790_ = _0788_ & ~(_0789_);
  assign _0791_ = _0790_ ^ _0787_;
  assign _0792_ = ~(b_i[3] & a_i[6]);
  assign _0793_ = ~(b_i[4] & a_i[5]);
  assign _0794_ = _0793_ ^ _0792_;
  assign _0795_ = ~(b_i[5] & a_i[4]);
  assign _0796_ = _0795_ ^ _0794_;
  assign _0797_ = _0796_ ^ _0791_;
  assign _0798_ = _0705_ | _0698_;
  assign _0799_ = _0706_ & ~(_0711_);
  assign _0800_ = _0798_ & ~(_0799_);
  assign _0801_ = _0800_ ^ _0797_;
  assign _0802_ = _0708_ | _0707_;
  assign _0803_ = _0709_ & ~(_0710_);
  assign _0804_ = _0802_ & ~(_0803_);
  assign _0805_ = ~(b_i[6] & a_i[3]);
  assign _0806_ = b_i[7] & a_i[2];
  assign _0807_ = ~(_0806_ ^ _0805_);
  assign _0808_ = b_i[8] & a_i[1];
  assign _0809_ = ~_0808_;
  assign _0810_ = _0809_ ^ _0807_;
  assign _0811_ = _0810_ ^ _0804_;
  assign _0812_ = _0730_ | ~(_0731_);
  assign _0813_ = _0732_ & ~(_0734_);
  assign _0814_ = _0812_ & ~(_0813_);
  assign _0815_ = _0814_ ^ _0811_;
  assign _0816_ = _0815_ ^ _0801_;
  assign _0817_ = _0725_ | _0712_;
  assign _0818_ = _0726_ & ~(_0741_);
  assign _0819_ = _0817_ & ~(_0818_);
  assign _0820_ = _0819_ ^ _0816_;
  assign _0821_ = ~(_0735_ | _0729_);
  assign _0822_ = _0736_ & ~(_0740_);
  assign _0823_ = ~(_0822_ | _0821_);
  assign _0824_ = b_i[9] & a_i[0];
  assign _0825_ = _0824_ ^ _0823_;
  assign _0826_ = _0825_ ^ _0820_;
  assign _0827_ = ~_0826_;
  assign _0828_ = _0755_ | _0742_;
  assign _0829_ = _0756_ & ~(_0758_);
  assign _0830_ = _0828_ & ~(_0829_);
  assign _0831_ = _0830_ ^ _0827_;
  assign _0832_ = _0760_ & ~(_0769_);
  assign _0833_ = _0832_ ^ _0831_;
  assign _0834_ = _0773_ & ~(_0770_);
  assign _0835_ = _0834_ ^ _0833_;
  assign _0836_ = _0777_ | _0774_;
  assign _0837_ = _0781_ & ~(_0778_);
  assign _0838_ = _0836_ & ~(_0837_);
  assign o[9] = _0838_ ^ _0835_;
  assign _0839_ = ~(a_i[10] & b_i[0]);
  assign _0840_ = ~(b_i[1] & a_i[9]);
  assign _0841_ = _0840_ ^ _0839_;
  assign _0842_ = ~(b_i[2] & a_i[8]);
  assign _0843_ = _0842_ ^ _0841_;
  assign _0844_ = _0784_ | _0783_;
  assign _0845_ = _0785_ & ~(_0786_);
  assign _0846_ = _0844_ & ~(_0845_);
  assign _0847_ = _0846_ ^ _0843_;
  assign _0848_ = ~(b_i[3] & a_i[7]);
  assign _0849_ = b_i[4] & a_i[6];
  assign _0850_ = ~(_0849_ ^ _0848_);
  assign _0851_ = b_i[5] & a_i[5];
  assign _0852_ = ~_0851_;
  assign _0853_ = _0852_ ^ _0850_;
  assign _0854_ = _0853_ ^ _0847_;
  assign _0855_ = _0790_ | _0787_;
  assign _0856_ = _0791_ & ~(_0796_);
  assign _0857_ = _0855_ & ~(_0856_);
  assign _0858_ = _0857_ ^ _0854_;
  assign _0859_ = _0793_ | _0792_;
  assign _0860_ = _0794_ & ~(_0795_);
  assign _0861_ = _0859_ & ~(_0860_);
  assign _0862_ = ~(b_i[6] & a_i[4]);
  assign _0863_ = b_i[7] & a_i[3];
  assign _0864_ = _0863_ ^ _0862_;
  assign _0865_ = b_i[8] & a_i[2];
  assign _0866_ = _0865_ ^ _0864_;
  assign _0867_ = _0866_ ^ _0861_;
  assign _0868_ = _0805_ | ~(_0806_);
  assign _0869_ = _0807_ & ~(_0809_);
  assign _0870_ = _0868_ & ~(_0869_);
  assign _0871_ = _0870_ ^ _0867_;
  assign _0872_ = _0871_ ^ _0858_;
  assign _0873_ = _0800_ | _0797_;
  assign _0874_ = _0801_ & ~(_0815_);
  assign _0875_ = _0873_ & ~(_0874_);
  assign _0876_ = _0875_ ^ _0872_;
  assign _0877_ = ~(_0810_ | _0804_);
  assign _0878_ = _0811_ & ~(_0814_);
  assign _0879_ = _0878_ | _0877_;
  assign _0880_ = b_i[9] & a_i[1];
  assign _0881_ = b_i[10] & a_i[0];
  assign _0882_ = ~(_0881_ ^ _0880_);
  assign _0883_ = _0882_ ^ _0879_;
  assign _0884_ = _0883_ ^ _0876_;
  assign _0885_ = _0819_ | _0816_;
  assign _0886_ = _0820_ & ~(_0825_);
  assign _0887_ = _0885_ & ~(_0886_);
  assign _0888_ = _0887_ ^ _0884_;
  assign _0889_ = _0824_ & ~(_0823_);
  assign _0890_ = ~_0889_;
  assign _0891_ = _0890_ ^ _0888_;
  assign _0892_ = _0827_ & ~(_0830_);
  assign _0893_ = _0892_ ^ _0891_;
  assign _0894_ = _0831_ | ~(_0832_);
  assign _0895_ = ~(_0894_ ^ _0893_);
  assign _0896_ = _0834_ & ~(_0833_);
  assign _0897_ = ~(_0836_ | _0835_);
  assign _0898_ = _0897_ | _0896_;
  assign _0899_ = _0835_ | _0778_;
  assign _0900_ = _0899_ | _0782_;
  assign _0901_ = _0900_ & ~(_0898_);
  assign o[10] = _0901_ ^ _0895_;
  assign _0902_ = ~(a_i[11] & b_i[0]);
  assign _0903_ = ~(b_i[1] & a_i[10]);
  assign _0904_ = _0903_ ^ _0902_;
  assign _0905_ = ~(b_i[2] & a_i[9]);
  assign _0906_ = _0905_ ^ _0904_;
  assign _0907_ = _0840_ | _0839_;
  assign _0908_ = _0841_ & ~(_0842_);
  assign _0909_ = _0907_ & ~(_0908_);
  assign _0910_ = _0909_ ^ _0906_;
  assign _0911_ = ~(b_i[3] & a_i[8]);
  assign _0912_ = ~(b_i[4] & a_i[7]);
  assign _0913_ = _0912_ ^ _0911_;
  assign _0914_ = ~(b_i[5] & a_i[6]);
  assign _0915_ = _0914_ ^ _0913_;
  assign _0916_ = _0915_ ^ _0910_;
  assign _0917_ = _0846_ | _0843_;
  assign _0918_ = _0847_ & ~(_0853_);
  assign _0919_ = _0917_ & ~(_0918_);
  assign _0920_ = _0919_ ^ _0916_;
  assign _0921_ = _0848_ | ~(_0849_);
  assign _0922_ = _0850_ & ~(_0852_);
  assign _0923_ = _0921_ & ~(_0922_);
  assign _0924_ = ~(b_i[6] & a_i[5]);
  assign _0925_ = ~(b_i[7] & a_i[4]);
  assign _0926_ = _0925_ ^ _0924_;
  assign _0927_ = ~(b_i[8] & a_i[3]);
  assign _0928_ = _0927_ ^ _0926_;
  assign _0929_ = _0928_ ^ _0923_;
  assign _0930_ = _0862_ | ~(_0863_);
  assign _0931_ = _0865_ & ~(_0864_);
  assign _0932_ = _0930_ & ~(_0931_);
  assign _0933_ = _0932_ ^ _0929_;
  assign _0934_ = _0933_ ^ _0920_;
  assign _0935_ = _0857_ | _0854_;
  assign _0936_ = _0858_ & ~(_0871_);
  assign _0937_ = _0935_ & ~(_0936_);
  assign _0938_ = _0937_ ^ _0934_;
  assign _0939_ = ~(_0866_ | _0861_);
  assign _0940_ = _0867_ & ~(_0870_);
  assign _0941_ = _0940_ | _0939_;
  assign _0942_ = ~(b_i[9] & a_i[2]);
  assign _0943_ = ~(b_i[10] & a_i[1]);
  assign _0944_ = _0943_ ^ _0942_;
  assign _0945_ = ~(b_i[11] & a_i[0]);
  assign _0946_ = _0945_ ^ _0944_;
  assign _0947_ = _0881_ & _0880_;
  assign _0948_ = _0947_ ^ _0946_;
  assign _0949_ = _0948_ ^ _0941_;
  assign _0950_ = _0949_ ^ _0938_;
  assign _0951_ = _0875_ | _0872_;
  assign _0952_ = _0876_ & ~(_0883_);
  assign _0953_ = _0951_ & ~(_0952_);
  assign _0954_ = _0953_ ^ _0950_;
  assign _0955_ = _0879_ & ~(_0882_);
  assign _0956_ = ~_0955_;
  assign _0957_ = _0956_ ^ _0954_;
  assign _0958_ = _0887_ | _0884_;
  assign _0959_ = _0888_ & ~(_0890_);
  assign _0960_ = _0958_ & ~(_0959_);
  assign _0961_ = _0960_ ^ _0957_;
  assign _0962_ = _0891_ | ~(_0892_);
  assign _0963_ = _0962_ ^ _0961_;
  assign _0964_ = _0894_ | _0893_;
  assign _0965_ = ~(_0901_ | _0895_);
  assign _0966_ = _0964_ & ~(_0965_);
  assign o[11] = _0966_ ^ _0963_;
  assign _0967_ = ~(a_i[12] & b_i[0]);
  assign _0968_ = ~(b_i[1] & a_i[11]);
  assign _0969_ = _0968_ ^ _0967_;
  assign _0970_ = ~(b_i[2] & a_i[10]);
  assign _0971_ = _0970_ ^ _0969_;
  assign _0972_ = _0903_ | _0902_;
  assign _0973_ = _0904_ & ~(_0905_);
  assign _0974_ = _0972_ & ~(_0973_);
  assign _0975_ = _0974_ ^ _0971_;
  assign _0976_ = ~(b_i[3] & a_i[9]);
  assign _0977_ = ~(b_i[4] & a_i[8]);
  assign _0978_ = _0977_ ^ _0976_;
  assign _0979_ = ~(b_i[5] & a_i[7]);
  assign _0980_ = _0979_ ^ _0978_;
  assign _0981_ = _0980_ ^ _0975_;
  assign _0982_ = _0909_ | _0906_;
  assign _0983_ = _0910_ & ~(_0915_);
  assign _0984_ = _0982_ & ~(_0983_);
  assign _0985_ = _0984_ ^ _0981_;
  assign _0986_ = _0912_ | _0911_;
  assign _0987_ = _0913_ & ~(_0914_);
  assign _0988_ = _0986_ & ~(_0987_);
  assign _0989_ = ~(b_i[6] & a_i[6]);
  assign _0990_ = ~(b_i[7] & a_i[5]);
  assign _0991_ = _0990_ ^ _0989_;
  assign _0992_ = ~(b_i[8] & a_i[4]);
  assign _0993_ = _0992_ ^ _0991_;
  assign _0994_ = _0993_ ^ _0988_;
  assign _0995_ = _0925_ | _0924_;
  assign _0996_ = _0926_ & ~(_0927_);
  assign _0997_ = _0995_ & ~(_0996_);
  assign _0998_ = _0997_ ^ _0994_;
  assign _0999_ = _0998_ ^ _0985_;
  assign _1000_ = _0919_ | _0916_;
  assign _1001_ = _0920_ & ~(_0933_);
  assign _1002_ = _1000_ & ~(_1001_);
  assign _1003_ = _1002_ ^ _0999_;
  assign _1004_ = _0928_ | _0923_;
  assign _1005_ = _0929_ & ~(_0932_);
  assign _1006_ = _1004_ & ~(_1005_);
  assign _1007_ = ~(b_i[9] & a_i[3]);
  assign _1008_ = ~(b_i[10] & a_i[2]);
  assign _1009_ = _1008_ ^ _1007_;
  assign _1010_ = ~(b_i[11] & a_i[1]);
  assign _1011_ = _1010_ ^ _1009_;
  assign _1012_ = _0943_ | _0942_;
  assign _1013_ = _0944_ & ~(_0945_);
  assign _1014_ = _1012_ & ~(_1013_);
  assign _1015_ = _1014_ ^ _1011_;
  assign _1016_ = b_i[12] & a_i[0];
  assign _1017_ = ~_1016_;
  assign _1018_ = _1017_ ^ _1015_;
  assign _1019_ = ~(_1018_ ^ _1006_);
  assign _1020_ = _0947_ & ~(_0946_);
  assign _1021_ = _1020_ ^ _1019_;
  assign _1022_ = _1021_ ^ _1003_;
  assign _1023_ = _0937_ | _0934_;
  assign _1024_ = _0938_ & ~(_0949_);
  assign _1025_ = _1023_ & ~(_1024_);
  assign _1026_ = _1025_ ^ _1022_;
  assign _1027_ = _0941_ & ~(_0948_);
  assign _1028_ = _1027_ ^ _1026_;
  assign _1029_ = _0953_ | _0950_;
  assign _1030_ = _0954_ & ~(_0956_);
  assign _1031_ = _1029_ & ~(_1030_);
  assign _1032_ = _1031_ ^ _1028_;
  assign _1033_ = _0960_ | _0957_;
  assign _1034_ = ~(_1033_ ^ _1032_);
  assign _1035_ = _0961_ & ~(_0962_);
  assign _1036_ = ~(_0964_ | _0963_);
  assign _1037_ = _1036_ | _1035_;
  assign _1038_ = _0963_ | _0895_;
  assign _1039_ = _0898_ & ~(_1038_);
  assign _1040_ = _1039_ | _1037_;
  assign _1041_ = _1038_ | _0899_;
  assign _1042_ = _0781_ & ~(_1041_);
  assign _1043_ = ~(_1042_ | _1040_);
  assign o[12] = _1043_ ^ _1034_;
  assign _1044_ = ~(a_i[13] & b_i[0]);
  assign _1045_ = ~(b_i[1] & a_i[12]);
  assign _1046_ = _1045_ ^ _1044_;
  assign _1047_ = ~(b_i[2] & a_i[11]);
  assign _1048_ = _1047_ ^ _1046_;
  assign _1049_ = _0968_ | _0967_;
  assign _1050_ = _0969_ & ~(_0970_);
  assign _1051_ = _1049_ & ~(_1050_);
  assign _1052_ = _1051_ ^ _1048_;
  assign _1053_ = ~(b_i[3] & a_i[10]);
  assign _1054_ = ~(b_i[4] & a_i[9]);
  assign _1055_ = _1054_ ^ _1053_;
  assign _1056_ = ~(b_i[5] & a_i[8]);
  assign _1057_ = _1056_ ^ _1055_;
  assign _1058_ = _1057_ ^ _1052_;
  assign _1059_ = _0974_ | _0971_;
  assign _1060_ = _0975_ & ~(_0980_);
  assign _1061_ = _1059_ & ~(_1060_);
  assign _1062_ = _1061_ ^ _1058_;
  assign _1063_ = _0977_ | _0976_;
  assign _1064_ = _0978_ & ~(_0979_);
  assign _1065_ = _1063_ & ~(_1064_);
  assign _1066_ = ~(b_i[6] & a_i[7]);
  assign _1067_ = b_i[7] & a_i[6];
  assign _1068_ = ~(_1067_ ^ _1066_);
  assign _1069_ = b_i[8] & a_i[5];
  assign _1070_ = ~_1069_;
  assign _1071_ = _1070_ ^ _1068_;
  assign _1072_ = _1071_ ^ _1065_;
  assign _1073_ = _0990_ | _0989_;
  assign _1074_ = _0991_ & ~(_0992_);
  assign _1075_ = _1073_ & ~(_1074_);
  assign _1076_ = _1075_ ^ _1072_;
  assign _1077_ = _1076_ ^ _1062_;
  assign _1078_ = _0984_ | _0981_;
  assign _1079_ = _0985_ & ~(_0998_);
  assign _1080_ = _1078_ & ~(_1079_);
  assign _1081_ = _1080_ ^ _1077_;
  assign _1082_ = _0993_ | _0988_;
  assign _1083_ = _0994_ & ~(_0997_);
  assign _1084_ = _1082_ & ~(_1083_);
  assign _1085_ = ~(b_i[9] & a_i[4]);
  assign _1086_ = ~(b_i[10] & a_i[3]);
  assign _1087_ = _1086_ ^ _1085_;
  assign _1088_ = ~(b_i[11] & a_i[2]);
  assign _1089_ = _1088_ ^ _1087_;
  assign _1090_ = _1008_ | _1007_;
  assign _1091_ = _1009_ & ~(_1010_);
  assign _1092_ = _1090_ & ~(_1091_);
  assign _1093_ = _1092_ ^ _1089_;
  assign _1094_ = b_i[12] & a_i[1];
  assign _1095_ = b_i[13] & a_i[0];
  assign _1096_ = ~(_1095_ ^ _1094_);
  assign _1097_ = _1096_ ^ _1093_;
  assign _1098_ = _1097_ ^ _1084_;
  assign _1099_ = _1014_ | _1011_;
  assign _1100_ = _1015_ & ~(_1017_);
  assign _1101_ = _1099_ & ~(_1100_);
  assign _1102_ = _1101_ ^ _1098_;
  assign _1103_ = _1102_ ^ _1081_;
  assign _1104_ = _1002_ | _0999_;
  assign _1105_ = _1003_ & ~(_1021_);
  assign _1106_ = _1104_ & ~(_1105_);
  assign _1107_ = _1106_ ^ _1103_;
  assign _1108_ = _1018_ | _1006_;
  assign _1109_ = _1020_ & ~(_1019_);
  assign _1110_ = _1108_ & ~(_1109_);
  assign _1111_ = _1110_ ^ _1107_;
  assign _1112_ = _1025_ | _1022_;
  assign _1113_ = _1027_ & _1026_;
  assign _1114_ = _1112_ & ~(_1113_);
  assign _1115_ = ~(_1114_ ^ _1111_);
  assign _1116_ = _1028_ & ~(_1031_);
  assign _1117_ = _1116_ ^ _1115_;
  assign _1118_ = _1033_ | _1032_;
  assign _1119_ = ~(_1043_ | _1034_);
  assign _1120_ = _1118_ & ~(_1119_);
  assign o[13] = _1120_ ^ _1117_;
  assign _1121_ = ~(a_i[14] & b_i[0]);
  assign _1122_ = ~(b_i[1] & a_i[13]);
  assign _1123_ = _1122_ ^ _1121_;
  assign _1124_ = ~(b_i[2] & a_i[12]);
  assign _1125_ = _1124_ ^ _1123_;
  assign _1126_ = _1045_ | _1044_;
  assign _1127_ = _1046_ & ~(_1047_);
  assign _1128_ = _1126_ & ~(_1127_);
  assign _1129_ = _1128_ ^ _1125_;
  assign _1130_ = ~(b_i[3] & a_i[11]);
  assign _1131_ = ~(b_i[4] & a_i[10]);
  assign _1132_ = _1131_ ^ _1130_;
  assign _1133_ = ~(b_i[5] & a_i[9]);
  assign _1134_ = _1133_ ^ _1132_;
  assign _1135_ = _1134_ ^ _1129_;
  assign _1136_ = _1051_ | _1048_;
  assign _1137_ = _1052_ & ~(_1057_);
  assign _1138_ = _1136_ & ~(_1137_);
  assign _1139_ = _1138_ ^ _1135_;
  assign _1140_ = _1054_ | _1053_;
  assign _1141_ = _1055_ & ~(_1056_);
  assign _1142_ = _1140_ & ~(_1141_);
  assign _1143_ = ~(b_i[6] & a_i[8]);
  assign _1144_ = b_i[7] & a_i[7];
  assign _1145_ = ~(_1144_ ^ _1143_);
  assign _1146_ = b_i[8] & a_i[6];
  assign _1147_ = ~_1146_;
  assign _1148_ = _1147_ ^ _1145_;
  assign _1149_ = _1148_ ^ _1142_;
  assign _1150_ = _1066_ | ~(_1067_);
  assign _1151_ = _1068_ & ~(_1070_);
  assign _1152_ = _1150_ & ~(_1151_);
  assign _1153_ = _1152_ ^ _1149_;
  assign _1154_ = _1153_ ^ _1139_;
  assign _1155_ = _1061_ | _1058_;
  assign _1156_ = _1062_ & ~(_1076_);
  assign _1157_ = _1155_ & ~(_1156_);
  assign _1158_ = _1157_ ^ _1154_;
  assign _1159_ = _1071_ | _1065_;
  assign _1160_ = _1072_ & ~(_1075_);
  assign _1161_ = _1159_ & ~(_1160_);
  assign _1162_ = ~(b_i[9] & a_i[5]);
  assign _1163_ = b_i[10] & a_i[4];
  assign _1164_ = ~(_1163_ ^ _1162_);
  assign _1165_ = b_i[11] & a_i[3];
  assign _1166_ = ~_1165_;
  assign _1167_ = _1166_ ^ _1164_;
  assign _1168_ = _1086_ | _1085_;
  assign _1169_ = _1087_ & ~(_1088_);
  assign _1170_ = _1168_ & ~(_1169_);
  assign _1171_ = _1170_ ^ _1167_;
  assign _1172_ = b_i[12] & a_i[2];
  assign _1173_ = b_i[13] & a_i[1];
  assign _1174_ = ~(_1173_ ^ _1172_);
  assign _1175_ = b_i[14] & a_i[0];
  assign _1176_ = _1175_ ^ _1174_;
  assign _1177_ = _1176_ ^ _1171_;
  assign _1178_ = _1177_ ^ _1161_;
  assign _1179_ = _1092_ | _1089_;
  assign _1180_ = _1093_ & ~(_1096_);
  assign _1181_ = _1179_ & ~(_1180_);
  assign _1182_ = _1181_ ^ _1178_;
  assign _1183_ = _1182_ ^ _1158_;
  assign _1184_ = _1080_ | _1077_;
  assign _1185_ = _1081_ & ~(_1102_);
  assign _1186_ = _1184_ & ~(_1185_);
  assign _1187_ = _1186_ ^ _1183_;
  assign _1188_ = _1097_ | _1084_;
  assign _1190_ = _1098_ & ~(_1101_);
  assign _1191_ = _1188_ & ~(_1190_);
  assign _1192_ = _1095_ & _1094_;
  assign _1193_ = _1192_ ^ _1191_;
  assign _1194_ = ~(_1193_ ^ _1187_);
  assign _1195_ = _1106_ | _1103_;
  assign _1196_ = _1107_ & ~(_1110_);
  assign _1197_ = _1195_ & ~(_1196_);
  assign _1198_ = _1197_ ^ _1194_;
  assign _1199_ = _1114_ | _1111_;
  assign _1201_ = ~(_1199_ ^ _1198_);
  assign _1202_ = _1116_ & ~(_1115_);
  assign _1203_ = ~(_1118_ | _1117_);
  assign _1204_ = _1203_ | _1202_;
  assign _1205_ = _1117_ | _1034_;
  assign _1206_ = _1205_ | _1043_;
  assign _1207_ = _1206_ & ~(_1204_);
  assign o[14] = _1207_ ^ _1201_;
  assign _1208_ = ~(a_i[15] & b_i[0]);
  assign _1209_ = ~(b_i[1] & a_i[14]);
  assign _1211_ = _1209_ ^ _1208_;
  assign _1212_ = ~(b_i[2] & a_i[13]);
  assign _1213_ = _1212_ ^ _1211_;
  assign _1214_ = _1122_ | _1121_;
  assign _1215_ = _1123_ & ~(_1124_);
  assign _1216_ = _1214_ & ~(_1215_);
  assign _1217_ = _1216_ ^ _1213_;
  assign _1218_ = ~(b_i[3] & a_i[12]);
  assign _1219_ = ~(b_i[4] & a_i[11]);
  assign _1220_ = _1219_ ^ _1218_;
  assign _1222_ = ~(b_i[5] & a_i[10]);
  assign _1223_ = _1222_ ^ _1220_;
  assign _1224_ = _1223_ ^ _1217_;
  assign _1225_ = _1128_ | _1125_;
  assign _1226_ = _1129_ & ~(_1134_);
  assign _1227_ = _1225_ & ~(_1226_);
  assign _1228_ = _1227_ ^ _1224_;
  assign _1229_ = _1131_ | _1130_;
  assign _1230_ = _1132_ & ~(_1133_);
  assign _1231_ = _1229_ & ~(_1230_);
  assign _1233_ = ~(b_i[6] & a_i[9]);
  assign _1234_ = b_i[7] & a_i[8];
  assign _1235_ = ~(_1234_ ^ _1233_);
  assign _1236_ = b_i[8] & a_i[7];
  assign _1237_ = ~_1236_;
  assign _1238_ = _1237_ ^ _1235_;
  assign _1239_ = _1238_ ^ _1231_;
  assign _1240_ = _1143_ | ~(_1144_);
  assign _1241_ = _1145_ & ~(_1147_);
  assign _1242_ = _1240_ & ~(_1241_);
  assign _1244_ = _1242_ ^ _1239_;
  assign _1245_ = _1244_ ^ _1228_;
  assign _1246_ = _1138_ | _1135_;
  assign _1247_ = _1139_ & ~(_1153_);
  assign _1248_ = _1246_ & ~(_1247_);
  assign _1249_ = _1248_ ^ _1245_;
  assign _1250_ = _1148_ | _1142_;
  assign _1251_ = _1149_ & ~(_1152_);
  assign _1252_ = _1250_ & ~(_1251_);
  assign _1253_ = b_i[9] & a_i[6];
  assign _1255_ = b_i[10] & a_i[5];
  assign _1256_ = _1255_ ^ _1253_;
  assign _1257_ = b_i[11] & a_i[4];
  assign _1258_ = ~_1257_;
  assign _1259_ = _1258_ ^ _1256_;
  assign _1260_ = _1162_ | ~(_1163_);
  assign _1261_ = _1164_ & ~(_1166_);
  assign _1262_ = _1260_ & ~(_1261_);
  assign _1263_ = _1262_ ^ _1259_;
  assign _1264_ = b_i[12] & a_i[3];
  assign _1266_ = b_i[13] & a_i[2];
  assign _1267_ = ~(_1266_ ^ _1264_);
  assign _1268_ = b_i[14] & a_i[1];
  assign _1269_ = _1268_ ^ _1267_;
  assign _1270_ = _1269_ ^ _1263_;
  assign _1271_ = _1270_ ^ _1252_;
  assign _1272_ = _1170_ | _1167_;
  assign _1273_ = _1171_ & ~(_1176_);
  assign _1274_ = _1272_ & ~(_1273_);
  assign _1275_ = _1274_ ^ _1271_;
  assign _1276_ = _1275_ ^ _1249_;
  assign _1277_ = _1157_ | _1154_;
  assign _1278_ = _1158_ & ~(_1182_);
  assign _1279_ = _1277_ & ~(_1278_);
  assign _1280_ = _1279_ ^ _1276_;
  assign _1281_ = _1177_ | _1161_;
  assign _1282_ = _1178_ & ~(_1181_);
  assign _1283_ = _1281_ & ~(_1282_);
  assign _1284_ = ~(_1173_ & _1172_);
  assign _1285_ = _1175_ & ~(_1174_);
  assign _1287_ = _1284_ & ~(_1285_);
  assign _1288_ = _1287_ ^ _1283_;
  assign _1289_ = b_i[15] & a_i[0];
  assign _1290_ = ~_1289_;
  assign _1291_ = _1290_ ^ _1288_;
  assign _1292_ = _1291_ ^ _1280_;
  assign _1293_ = _1186_ | _1183_;
  assign _1294_ = _1187_ & ~(_1193_);
  assign _1295_ = _1293_ & ~(_1294_);
  assign _1296_ = _1295_ ^ _1292_;
  assign _1298_ = _1192_ & ~(_1191_);
  assign _1299_ = _1298_ ^ _1296_;
  assign _1300_ = _1197_ | ~(_1194_);
  assign _1301_ = _1300_ ^ _1299_;
  assign _1302_ = _1199_ | _1198_;
  assign _1303_ = ~(_1207_ | _1201_);
  assign _1304_ = _1302_ & ~(_1303_);
  assign o[15] = _1304_ ^ _1301_;
  assign _1305_ = ~(b_i[1] & a_i[15]);
  assign _1306_ = b_i[2] & a_i[14];
  assign _1308_ = _1306_ ^ _1305_;
  assign _1309_ = _1209_ | _1208_;
  assign _1310_ = _1211_ & ~(_1212_);
  assign _1311_ = _1309_ & ~(_1310_);
  assign _1312_ = _1311_ ^ _1308_;
  assign _1313_ = ~(b_i[3] & a_i[13]);
  assign _1314_ = ~(b_i[4] & a_i[12]);
  assign _1315_ = _1314_ ^ _1313_;
  assign _1316_ = ~(b_i[5] & a_i[11]);
  assign _1317_ = _1316_ ^ _1315_;
  assign _1319_ = _1317_ ^ _1312_;
  assign _1320_ = _1216_ | _1213_;
  assign _1321_ = _1217_ & ~(_1223_);
  assign _1322_ = _1320_ & ~(_1321_);
  assign _1323_ = _1322_ ^ _1319_;
  assign _1324_ = _1219_ | _1218_;
  assign _1325_ = _1220_ & ~(_1222_);
  assign _1326_ = _1324_ & ~(_1325_);
  assign _1327_ = ~(b_i[6] & a_i[10]);
  assign _1328_ = b_i[7] & a_i[9];
  assign _1330_ = ~(_1328_ ^ _1327_);
  assign _1331_ = b_i[8] & a_i[8];
  assign _1332_ = ~_1331_;
  assign _1333_ = _1332_ ^ _1330_;
  assign _1334_ = _1333_ ^ _1326_;
  assign _1335_ = _1233_ | ~(_1234_);
  assign _1336_ = _1235_ & ~(_1237_);
  assign _1337_ = _1335_ & ~(_1336_);
  assign _1338_ = _1337_ ^ _1334_;
  assign _1339_ = _1338_ ^ _1323_;
  assign _1341_ = _1227_ | _1224_;
  assign _1342_ = _1228_ & ~(_1244_);
  assign _1343_ = _1341_ & ~(_1342_);
  assign _1344_ = _1343_ ^ _1339_;
  assign _1345_ = _1238_ | _1231_;
  assign _1346_ = _1239_ & ~(_1242_);
  assign _1347_ = _1345_ & ~(_1346_);
  assign _1348_ = b_i[9] & a_i[7];
  assign _1349_ = b_i[10] & a_i[6];
  assign _1350_ = _1349_ ^ _1348_;
  assign _1352_ = b_i[11] & a_i[5];
  assign _1353_ = ~_1352_;
  assign _1354_ = _1353_ ^ _1350_;
  assign _1355_ = ~(_1255_ & _1253_);
  assign _1356_ = _1256_ & ~(_1258_);
  assign _1357_ = _1355_ & ~(_1356_);
  assign _1358_ = _1357_ ^ _1354_;
  assign _1359_ = b_i[12] & a_i[4];
  assign _1360_ = b_i[13] & a_i[3];
  assign _1361_ = ~(_1360_ ^ _1359_);
  assign _1363_ = b_i[14] & a_i[2];
  assign _1364_ = _1363_ ^ _1361_;
  assign _1365_ = _1364_ ^ _1358_;
  assign _1366_ = _1365_ ^ _1347_;
  assign _1367_ = _1262_ | _1259_;
  assign _1368_ = _1263_ & ~(_1269_);
  assign _1369_ = _1367_ & ~(_1368_);
  assign _1370_ = _1369_ ^ _1366_;
  assign _1371_ = _1370_ ^ _1344_;
  assign _1372_ = _1248_ | _1245_;
  assign _1374_ = _1249_ & ~(_1275_);
  assign _1375_ = _1372_ & ~(_1374_);
  assign _1376_ = _1375_ ^ _1371_;
  assign _1377_ = _1270_ | _1252_;
  assign _1378_ = _1271_ & ~(_1274_);
  assign _1379_ = _1377_ & ~(_1378_);
  assign _1380_ = ~(_1266_ & _1264_);
  assign _1381_ = _1268_ & ~(_1267_);
  assign _1382_ = _1380_ & ~(_1381_);
  assign _1383_ = ~(_1382_ ^ _1379_);
  assign _1385_ = b_i[15] & a_i[1];
  assign _1386_ = _1385_ ^ _1383_;
  assign _1387_ = _1386_ ^ _1376_;
  assign _1388_ = _1279_ | _1276_;
  assign _1389_ = _1280_ & ~(_1291_);
  assign _1390_ = _1388_ & ~(_1389_);
  assign _1391_ = _1390_ ^ _1387_;
  assign _1392_ = _1287_ | _1283_;
  assign _1393_ = _1288_ & ~(_1290_);
  assign _1394_ = _1392_ & ~(_1393_);
  assign _1396_ = _1394_ ^ _1391_;
  assign _1397_ = _1295_ | _1292_;
  assign _1398_ = _1298_ & _1296_;
  assign _1399_ = _1397_ & ~(_1398_);
  assign _1400_ = ~(_1399_ ^ _1396_);
  assign _1401_ = _1299_ & ~(_1300_);
  assign _1402_ = ~(_1302_ | _1301_);
  assign _1403_ = _1402_ | _1401_;
  assign _1404_ = _1301_ | _1201_;
  assign _1405_ = _1204_ & ~(_1404_);
  assign _1407_ = _1405_ | _1403_;
  assign _1408_ = _1404_ | _1205_;
  assign _1409_ = _1040_ & ~(_1408_);
  assign _1410_ = _1409_ | _1407_;
  assign _1411_ = _1408_ | _1041_;
  assign _1412_ = _0781_ & ~(_1411_);
  assign _1413_ = _1412_ | _1410_;
  assign o[16] = ~(_1413_ ^ _1400_);
  assign _1414_ = b_i[2] & a_i[15];
  assign _1415_ = _1306_ & ~(_1305_);
  assign _1417_ = _1415_ ^ _1414_;
  assign _1418_ = ~(b_i[3] & a_i[14]);
  assign _1419_ = b_i[4] & a_i[13];
  assign _1420_ = ~(_1419_ ^ _1418_);
  assign _1421_ = b_i[5] & a_i[12];
  assign _1422_ = ~_1421_;
  assign _1423_ = _1422_ ^ _1420_;
  assign _1424_ = _1423_ ^ _1417_;
  assign _1425_ = _1311_ | _1308_;
  assign _1426_ = _1312_ & ~(_1317_);
  assign _1427_ = _1425_ & ~(_1426_);
  assign _1428_ = _1427_ ^ _1424_;
  assign _1429_ = _1314_ | _1313_;
  assign _1430_ = _1315_ & ~(_1316_);
  assign _1431_ = _1429_ & ~(_1430_);
  assign _1432_ = ~(b_i[6] & a_i[11]);
  assign _1433_ = b_i[7] & a_i[10];
  assign _1434_ = _1433_ ^ _1432_;
  assign _1435_ = b_i[8] & a_i[9];
  assign _1436_ = _1435_ ^ _1434_;
  assign _1438_ = _1436_ ^ _1431_;
  assign _1439_ = _1327_ | ~(_1328_);
  assign _1440_ = _1330_ & ~(_1332_);
  assign _1441_ = _1439_ & ~(_1440_);
  assign _1442_ = _1441_ ^ _1438_;
  assign _1443_ = _1442_ ^ _1428_;
  assign _1444_ = _1322_ | _1319_;
  assign _1445_ = _1323_ & ~(_1338_);
  assign _1446_ = _1444_ & ~(_1445_);
  assign _1447_ = _1446_ ^ _1443_;
  assign _1449_ = _1333_ | _1326_;
  assign _1450_ = _1334_ & ~(_1337_);
  assign _1451_ = _1449_ & ~(_1450_);
  assign _1452_ = b_i[9] & a_i[8];
  assign _1453_ = b_i[10] & a_i[7];
  assign _1454_ = _1453_ ^ _1452_;
  assign _1455_ = b_i[11] & a_i[6];
  assign _1456_ = ~_1455_;
  assign _1457_ = _1456_ ^ _1454_;
  assign _1458_ = ~(_1349_ & _1348_);
  assign _1460_ = _1350_ & ~(_1353_);
  assign _1461_ = _1458_ & ~(_1460_);
  assign _1462_ = _1461_ ^ _1457_;
  assign _1463_ = b_i[12] & a_i[5];
  assign _1464_ = b_i[13] & a_i[4];
  assign _1465_ = ~(_1464_ ^ _1463_);
  assign _1466_ = b_i[14] & a_i[3];
  assign _1467_ = _1466_ ^ _1465_;
  assign _1468_ = _1467_ ^ _1462_;
  assign _1469_ = _1468_ ^ _1451_;
  assign _1471_ = _1357_ | _1354_;
  assign _1472_ = _1358_ & ~(_1364_);
  assign _1473_ = _1471_ & ~(_1472_);
  assign _1474_ = _1473_ ^ _1469_;
  assign _1475_ = _1474_ ^ _1447_;
  assign _1476_ = _1343_ | _1339_;
  assign _1477_ = _1344_ & ~(_1370_);
  assign _1478_ = _1476_ & ~(_1477_);
  assign _1479_ = _1478_ ^ _1475_;
  assign _1480_ = _1365_ | _1347_;
  assign _1482_ = _1366_ & ~(_1369_);
  assign _1483_ = _1480_ & ~(_1482_);
  assign _1484_ = ~(_1360_ & _1359_);
  assign _1485_ = _1363_ & ~(_1361_);
  assign _1486_ = _1484_ & ~(_1485_);
  assign _1487_ = ~(_1486_ ^ _1483_);
  assign _1488_ = b_i[15] & a_i[2];
  assign _1489_ = _1488_ ^ _1487_;
  assign _1490_ = _1489_ ^ _1479_;
  assign _1491_ = _1375_ | _1371_;
  assign _1493_ = _1376_ & ~(_1386_);
  assign _1494_ = _1491_ & ~(_1493_);
  assign _1495_ = _1494_ ^ _1490_;
  assign _1496_ = _1382_ | _1379_;
  assign _1497_ = _1385_ & ~(_1383_);
  assign _1498_ = _1496_ & ~(_1497_);
  assign _1499_ = ~(_1498_ ^ _1495_);
  assign _1500_ = _1390_ | _1387_;
  assign _1501_ = _1391_ & ~(_1394_);
  assign _1502_ = _1500_ & ~(_1501_);
  assign _1504_ = _1502_ ^ _1499_;
  assign _1505_ = _1399_ | _1396_;
  assign _1506_ = _1413_ & ~(_1400_);
  assign _1507_ = _1505_ & ~(_1506_);
  assign o[17] = _1507_ ^ _1504_;
  assign _1508_ = b_i[3] & a_i[15];
  assign _1509_ = b_i[4] & a_i[14];
  assign _1510_ = _1509_ ^ _1508_;
  assign _1511_ = b_i[5] & a_i[13];
  assign _1512_ = ~_1511_;
  assign _1514_ = _1512_ ^ _1510_;
  assign _1515_ = ~(_1415_ & _1414_);
  assign _1516_ = _1417_ & ~(_1423_);
  assign _1517_ = _1515_ & ~(_1516_);
  assign _1518_ = _1517_ ^ _1514_;
  assign _1519_ = _1418_ | ~(_1419_);
  assign _1520_ = _1420_ & ~(_1422_);
  assign _1521_ = _1519_ & ~(_1520_);
  assign _1522_ = b_i[6] & a_i[12];
  assign _1523_ = b_i[7] & a_i[11];
  assign _1525_ = ~(_1523_ ^ _1522_);
  assign _1526_ = b_i[8] & a_i[10];
  assign _1527_ = _1526_ ^ _1525_;
  assign _1528_ = _1527_ ^ _1521_;
  assign _1529_ = _1432_ | ~(_1433_);
  assign _1530_ = _1435_ & ~(_1434_);
  assign _1531_ = _1529_ & ~(_1530_);
  assign _1532_ = _1531_ ^ _1528_;
  assign _1533_ = _1532_ ^ _1518_;
  assign _1534_ = _1427_ | _1424_;
  assign _1536_ = _1428_ & ~(_1442_);
  assign _1537_ = _1534_ & ~(_1536_);
  assign _1538_ = _1537_ ^ _1533_;
  assign _1539_ = _1436_ | _1431_;
  assign _1540_ = _1438_ & ~(_1441_);
  assign _1541_ = _1539_ & ~(_1540_);
  assign _1542_ = b_i[9] & a_i[9];
  assign _1543_ = b_i[10] & a_i[8];
  assign _1544_ = ~(_1543_ ^ _1542_);
  assign _1545_ = b_i[11] & a_i[7];
  assign _0000_ = _1545_ ^ _1544_;
  assign _0001_ = ~(_1453_ & _1452_);
  assign _0002_ = _1454_ & ~(_1456_);
  assign _0003_ = _0001_ & ~(_0002_);
  assign _0004_ = _0003_ ^ _0000_;
  assign _0005_ = b_i[12] & a_i[6];
  assign _0006_ = b_i[13] & a_i[5];
  assign _0007_ = ~(_0006_ ^ _0005_);
  assign _0008_ = b_i[14] & a_i[4];
  assign _0009_ = _0008_ ^ _0007_;
  assign _0011_ = _0009_ ^ _0004_;
  assign _0012_ = _0011_ ^ _1541_;
  assign _0013_ = _1461_ | _1457_;
  assign _0014_ = _1462_ & ~(_1467_);
  assign _0015_ = _0013_ & ~(_0014_);
  assign _0016_ = _0015_ ^ _0012_;
  assign _0017_ = _0016_ ^ _1538_;
  assign _0018_ = _1446_ | _1443_;
  assign _0019_ = _1447_ & ~(_1474_);
  assign _0020_ = _0018_ & ~(_0019_);
  assign _0022_ = _0020_ ^ _0017_;
  assign _0023_ = _1468_ | _1451_;
  assign _0024_ = _1469_ & ~(_1473_);
  assign _0025_ = _0023_ & ~(_0024_);
  assign _0026_ = ~(_1464_ & _1463_);
  assign _0027_ = _1466_ & ~(_1465_);
  assign _0028_ = _0026_ & ~(_0027_);
  assign _0029_ = ~(_0028_ ^ _0025_);
  assign _0030_ = b_i[15] & a_i[3];
  assign _0031_ = _0030_ ^ _0029_;
  assign _0033_ = _0031_ ^ _0022_;
  assign _0034_ = _1478_ | _1475_;
  assign _0035_ = _1479_ & ~(_1489_);
  assign _0036_ = _0034_ & ~(_0035_);
  assign _0037_ = _0036_ ^ _0033_;
  assign _0038_ = _1486_ | _1483_;
  assign _0039_ = _1488_ & ~(_1487_);
  assign _0040_ = _0038_ & ~(_0039_);
  assign _0041_ = _0040_ ^ _0037_;
  assign _0042_ = _1494_ | _1490_;
  assign _0044_ = _1495_ & ~(_1498_);
  assign _0045_ = _0042_ & ~(_0044_);
  assign _0046_ = ~(_0045_ ^ _0041_);
  assign _0047_ = _1499_ & ~(_1502_);
  assign _0048_ = ~(_1505_ | _1504_);
  assign _0049_ = _0048_ | _0047_;
  assign _0050_ = _1504_ | _1400_;
  assign _0051_ = _0050_ | ~(_1413_);
  assign _0052_ = _0051_ & ~(_0049_);
  assign o[18] = _0052_ ^ _0046_;
  assign _0054_ = b_i[4] & a_i[15];
  assign _0055_ = b_i[5] & a_i[14];
  assign _0056_ = ~(_0055_ ^ _0054_);
  assign _0057_ = ~_0056_;
  assign _0058_ = ~(_1509_ & _1508_);
  assign _0059_ = _1510_ & ~(_1512_);
  assign _0060_ = _0058_ & ~(_0059_);
  assign _0061_ = b_i[6] & a_i[13];
  assign _0062_ = b_i[7] & a_i[12];
  assign _0063_ = ~(_0062_ ^ _0061_);
  assign _0065_ = b_i[8] & a_i[11];
  assign _0066_ = _0065_ ^ _0063_;
  assign _0067_ = _0066_ ^ _0060_;
  assign _0068_ = ~(_1523_ & _1522_);
  assign _0069_ = _1526_ & ~(_1525_);
  assign _0070_ = _0068_ & ~(_0069_);
  assign _0071_ = _0070_ ^ _0067_;
  assign _0072_ = _0071_ ^ _0057_;
  assign _0073_ = _1517_ | _1514_;
  assign _0074_ = _1518_ & ~(_1532_);
  assign _0076_ = _0073_ & ~(_0074_);
  assign _0077_ = _0076_ ^ _0072_;
  assign _0078_ = _1527_ | _1521_;
  assign _0079_ = _1528_ & ~(_1531_);
  assign _0080_ = _0078_ & ~(_0079_);
  assign _0081_ = b_i[9] & a_i[10];
  assign _0082_ = b_i[10] & a_i[9];
  assign _0083_ = ~(_0082_ ^ _0081_);
  assign _0084_ = b_i[11] & a_i[8];
  assign _0085_ = _0084_ ^ _0083_;
  assign _0087_ = ~(_1543_ & _1542_);
  assign _0088_ = _1545_ & ~(_1544_);
  assign _0089_ = _0087_ & ~(_0088_);
  assign _0090_ = _0089_ ^ _0085_;
  assign _0091_ = b_i[12] & a_i[7];
  assign _0092_ = b_i[13] & a_i[6];
  assign _0093_ = ~(_0092_ ^ _0091_);
  assign _0094_ = b_i[14] & a_i[5];
  assign _0095_ = _0094_ ^ _0093_;
  assign _0096_ = _0095_ ^ _0090_;
  assign _0097_ = _0096_ ^ _0080_;
  assign _0098_ = _0003_ | _0000_;
  assign _0099_ = _0004_ & ~(_0009_);
  assign _0100_ = _0098_ & ~(_0099_);
  assign _0101_ = _0100_ ^ _0097_;
  assign _0102_ = _0101_ ^ _0077_;
  assign _0103_ = _1537_ | _1533_;
  assign _0104_ = _1538_ & ~(_0016_);
  assign _0105_ = _0103_ & ~(_0104_);
  assign _0106_ = _0105_ ^ _0102_;
  assign _0108_ = _0011_ | _1541_;
  assign _0109_ = _0012_ & ~(_0015_);
  assign _0110_ = _0108_ & ~(_0109_);
  assign _0111_ = ~(_0006_ & _0005_);
  assign _0112_ = _0008_ & ~(_0007_);
  assign _0113_ = _0111_ & ~(_0112_);
  assign _0114_ = ~(_0113_ ^ _0110_);
  assign _0115_ = b_i[15] & a_i[4];
  assign _0116_ = _0115_ ^ _0114_;
  assign _0117_ = _0116_ ^ _0106_;
  assign _0119_ = _0020_ | _0017_;
  assign _0120_ = _0022_ & ~(_0031_);
  assign _0121_ = _0119_ & ~(_0120_);
  assign _0122_ = _0121_ ^ _0117_;
  assign _0123_ = _0028_ | _0025_;
  assign _0124_ = _0030_ & ~(_0029_);
  assign _0125_ = _0123_ & ~(_0124_);
  assign _0126_ = ~(_0125_ ^ _0122_);
  assign _0127_ = _0036_ | _0033_;
  assign _0128_ = _0037_ & ~(_0040_);
  assign _0130_ = _0127_ & ~(_0128_);
  assign _0131_ = _0130_ ^ _0126_;
  assign _0132_ = _0045_ | _0041_;
  assign _0133_ = ~(_0052_ | _0046_);
  assign _0134_ = _0132_ & ~(_0133_);
  assign o[19] = _0134_ ^ _0131_;
  assign _0135_ = b_i[5] & a_i[15];
  assign _0136_ = ~(_0055_ & _0054_);
  assign _0137_ = b_i[6] & a_i[14];
  assign _0138_ = b_i[7] & a_i[13];
  assign _0140_ = ~(_0138_ ^ _0137_);
  assign _0141_ = b_i[8] & a_i[12];
  assign _0142_ = _0141_ ^ _0140_;
  assign _0143_ = _0142_ ^ _0136_;
  assign _0144_ = ~(_0062_ & _0061_);
  assign _0145_ = _0065_ & ~(_0063_);
  assign _0146_ = _0144_ & ~(_0145_);
  assign _0147_ = _0146_ ^ _0143_;
  assign _0148_ = _0147_ ^ _0135_;
  assign _0149_ = _0057_ & ~(_0071_);
  assign _0151_ = _0149_ ^ _0148_;
  assign _0152_ = ~_0151_;
  assign _0153_ = _0066_ | _0060_;
  assign _0154_ = _0067_ & ~(_0070_);
  assign _0155_ = _0153_ & ~(_0154_);
  assign _0156_ = b_i[9] & a_i[11];
  assign _0157_ = b_i[10] & a_i[10];
  assign _0158_ = ~(_0157_ ^ _0156_);
  assign _0159_ = b_i[11] & a_i[9];
  assign _0160_ = _0159_ ^ _0158_;
  assign _0162_ = ~(_0082_ & _0081_);
  assign _0163_ = _0084_ & ~(_0083_);
  assign _0164_ = _0162_ & ~(_0163_);
  assign _0165_ = _0164_ ^ _0160_;
  assign _0166_ = b_i[12] & a_i[8];
  assign _0167_ = b_i[13] & a_i[7];
  assign _0168_ = ~(_0167_ ^ _0166_);
  assign _0169_ = b_i[14] & a_i[6];
  assign _0170_ = _0169_ ^ _0168_;
  assign _0171_ = _0170_ ^ _0165_;
  assign _0173_ = _0171_ ^ _0155_;
  assign _0174_ = _0089_ | _0085_;
  assign _0175_ = _0090_ & ~(_0095_);
  assign _0176_ = _0174_ & ~(_0175_);
  assign _0177_ = _0176_ ^ _0173_;
  assign _0178_ = _0177_ ^ _0152_;
  assign _0179_ = _0076_ | _0072_;
  assign _0180_ = _0077_ & ~(_0101_);
  assign _0181_ = _0179_ & ~(_0180_);
  assign _0182_ = _0181_ ^ _0178_;
  assign _0184_ = _0096_ | _0080_;
  assign _0185_ = _0097_ & ~(_0100_);
  assign _0186_ = _0184_ & ~(_0185_);
  assign _0187_ = ~(_0092_ & _0091_);
  assign _0188_ = _0094_ & ~(_0093_);
  assign _0189_ = _0187_ & ~(_0188_);
  assign _0190_ = ~(_0189_ ^ _0186_);
  assign _0191_ = b_i[15] & a_i[5];
  assign _0192_ = _0191_ ^ _0190_;
  assign _0193_ = _0192_ ^ _0182_;
  assign _0195_ = _0105_ | _0102_;
  assign _0196_ = _0106_ & ~(_0116_);
  assign _0197_ = _0195_ & ~(_0196_);
  assign _0198_ = _0197_ ^ _0193_;
  assign _0199_ = _0113_ | _0110_;
  assign _0200_ = _0115_ & ~(_0114_);
  assign _0201_ = _0199_ & ~(_0200_);
  assign _0202_ = _0201_ ^ _0198_;
  assign _0203_ = _0121_ | _0117_;
  assign _0204_ = _0122_ & ~(_0125_);
  assign _0206_ = _0203_ & ~(_0204_);
  assign _0207_ = ~(_0206_ ^ _0202_);
  assign _0208_ = _0126_ & ~(_0130_);
  assign _0209_ = ~(_0132_ | _0131_);
  assign _0210_ = _0209_ | _0208_;
  assign _0211_ = _0131_ | _0046_;
  assign _0212_ = _0049_ & ~(_0211_);
  assign _0213_ = _0212_ | _0210_;
  assign _0214_ = _0211_ | _0050_;
  assign _0215_ = _1413_ & ~(_0214_);
  assign _0217_ = ~(_0215_ | _0213_);
  assign o[20] = _0217_ ^ _0207_;
  assign _0218_ = b_i[6] & a_i[15];
  assign _0219_ = b_i[7] & a_i[14];
  assign _0220_ = ~(_0219_ ^ _0218_);
  assign _0221_ = b_i[8] & a_i[13];
  assign _0222_ = _0221_ ^ _0220_;
  assign _0223_ = ~(_0138_ & _0137_);
  assign _0224_ = _0141_ & ~(_0140_);
  assign _0225_ = _0223_ & ~(_0224_);
  assign _0227_ = ~(_0225_ ^ _0222_);
  assign _0228_ = _0135_ & ~(_0147_);
  assign _0229_ = _0228_ ^ _0227_;
  assign _0230_ = ~_0229_;
  assign _0231_ = _0142_ | _0136_;
  assign _0232_ = _0143_ & ~(_0146_);
  assign _0233_ = _0231_ & ~(_0232_);
  assign _0234_ = b_i[9] & a_i[12];
  assign _0235_ = b_i[10] & a_i[11];
  assign _0236_ = ~(_0235_ ^ _0234_);
  assign _0238_ = b_i[11] & a_i[10];
  assign _0239_ = _0238_ ^ _0236_;
  assign _0240_ = ~(_0157_ & _0156_);
  assign _0241_ = _0159_ & ~(_0158_);
  assign _0242_ = _0240_ & ~(_0241_);
  assign _0243_ = _0242_ ^ _0239_;
  assign _0244_ = b_i[12] & a_i[9];
  assign _0245_ = b_i[13] & a_i[8];
  assign _0246_ = ~(_0245_ ^ _0244_);
  assign _0247_ = b_i[14] & a_i[7];
  assign _0249_ = _0247_ ^ _0246_;
  assign _0250_ = _0249_ ^ _0243_;
  assign _0251_ = _0250_ ^ _0233_;
  assign _0252_ = _0164_ | _0160_;
  assign _0253_ = _0165_ & ~(_0170_);
  assign _0254_ = _0252_ & ~(_0253_);
  assign _0255_ = _0254_ ^ _0251_;
  assign _0256_ = _0255_ ^ _0230_;
  assign _0257_ = _0148_ | ~(_0149_);
  assign _0258_ = _0152_ & ~(_0177_);
  assign _0260_ = _0257_ & ~(_0258_);
  assign _0261_ = _0260_ ^ _0256_;
  assign _0262_ = _0171_ | _0155_;
  assign _0263_ = _0173_ & ~(_0176_);
  assign _0264_ = _0262_ & ~(_0263_);
  assign _0265_ = ~(_0167_ & _0166_);
  assign _0266_ = _0169_ & ~(_0168_);
  assign _0267_ = _0265_ & ~(_0266_);
  assign _0268_ = ~(_0267_ ^ _0264_);
  assign _0269_ = b_i[15] & a_i[6];
  assign _0271_ = _0269_ ^ _0268_;
  assign _0272_ = _0271_ ^ _0261_;
  assign _0273_ = _0181_ | _0178_;
  assign _0274_ = _0182_ & ~(_0192_);
  assign _0275_ = _0273_ & ~(_0274_);
  assign _0276_ = _0275_ ^ _0272_;
  assign _0277_ = _0189_ | _0186_;
  assign _0278_ = _0191_ & ~(_0190_);
  assign _0279_ = _0277_ & ~(_0278_);
  assign _0280_ = _0279_ ^ _0276_;
  assign _0282_ = ~_0280_;
  assign _0283_ = _0197_ | _0193_;
  assign _0284_ = _0198_ & ~(_0201_);
  assign _0285_ = _0283_ & ~(_0284_);
  assign _0286_ = _0285_ ^ _0282_;
  assign _0287_ = _0206_ | _0202_;
  assign _0288_ = ~(_0217_ | _0207_);
  assign _0289_ = _0287_ & ~(_0288_);
  assign o[21] = _0289_ ^ _0286_;
  assign _0290_ = b_i[7] & a_i[15];
  assign _0292_ = b_i[8] & a_i[14];
  assign _0293_ = ~(_0292_ ^ _0290_);
  assign _0294_ = ~(_0219_ & _0218_);
  assign _0295_ = _0221_ & ~(_0220_);
  assign _0296_ = _0294_ & ~(_0295_);
  assign _0297_ = ~(_0296_ ^ _0293_);
  assign _0298_ = ~_0297_;
  assign _0299_ = _0225_ | _0222_;
  assign _0300_ = b_i[9] & a_i[13];
  assign _0301_ = b_i[10] & a_i[12];
  assign _0303_ = ~(_0301_ ^ _0300_);
  assign _0304_ = b_i[11] & a_i[11];
  assign _0305_ = _0304_ ^ _0303_;
  assign _0306_ = ~(_0235_ & _0234_);
  assign _0307_ = _0238_ & ~(_0236_);
  assign _0308_ = _0306_ & ~(_0307_);
  assign _0309_ = _0308_ ^ _0305_;
  assign _0310_ = b_i[12] & a_i[10];
  assign _0311_ = b_i[13] & a_i[9];
  assign _0312_ = ~(_0311_ ^ _0310_);
  assign _0314_ = b_i[14] & a_i[8];
  assign _0315_ = _0314_ ^ _0312_;
  assign _0316_ = _0315_ ^ _0309_;
  assign _0317_ = _0316_ ^ _0299_;
  assign _0318_ = _0242_ | _0239_;
  assign _0319_ = _0243_ & ~(_0249_);
  assign _0320_ = _0318_ & ~(_0319_);
  assign _0321_ = _0320_ ^ _0317_;
  assign _0322_ = _0321_ ^ _0298_;
  assign _0323_ = _0227_ | ~(_0228_);
  assign _0325_ = _0230_ & ~(_0255_);
  assign _0326_ = _0323_ & ~(_0325_);
  assign _0327_ = ~(_0326_ ^ _0322_);
  assign _0328_ = _0250_ | _0233_;
  assign _0329_ = _0251_ & ~(_0254_);
  assign _0330_ = _0328_ & ~(_0329_);
  assign _0331_ = ~(_0245_ & _0244_);
  assign _0332_ = _0247_ & ~(_0246_);
  assign _0333_ = _0331_ & ~(_0332_);
  assign _0334_ = ~(_0333_ ^ _0330_);
  assign _0336_ = b_i[15] & a_i[7];
  assign _0337_ = _0336_ ^ _0334_;
  assign _0338_ = ~(_0337_ ^ _0327_);
  assign _0339_ = _0260_ | _0256_;
  assign _0340_ = _0261_ & ~(_0271_);
  assign _0341_ = _0339_ & ~(_0340_);
  assign _0342_ = _0341_ ^ _0338_;
  assign _0343_ = _0267_ | _0264_;
  assign _0344_ = _0269_ & ~(_0268_);
  assign _0345_ = _0343_ & ~(_0344_);
  assign _0347_ = _0345_ ^ _0342_;
  assign _0348_ = _0275_ | _0272_;
  assign _0349_ = _0276_ & ~(_0279_);
  assign _0350_ = _0348_ & ~(_0349_);
  assign _0351_ = ~(_0350_ ^ _0347_);
  assign _0352_ = _0282_ & ~(_0285_);
  assign _0353_ = ~(_0287_ | _0286_);
  assign _0354_ = _0353_ | _0352_;
  assign _0355_ = _0286_ | _0207_;
  assign _0356_ = _0355_ | _0217_;
  assign _0358_ = _0356_ & ~(_0354_);
  assign o[22] = _0358_ ^ _0351_;
  assign _0359_ = b_i[8] & a_i[15];
  assign _0360_ = ~_0359_;
  assign _0361_ = _0292_ & _0290_;
  assign _0362_ = _0361_ ^ _0360_;
  assign _0363_ = ~_0362_;
  assign _0364_ = _0296_ | _0293_;
  assign _0365_ = b_i[9] & a_i[14];
  assign _0366_ = b_i[10] & a_i[13];
  assign _0368_ = ~(_0366_ ^ _0365_);
  assign _0369_ = b_i[11] & a_i[12];
  assign _0370_ = _0369_ ^ _0368_;
  assign _0371_ = ~(_0301_ & _0300_);
  assign _0372_ = _0304_ & ~(_0303_);
  assign _0373_ = _0371_ & ~(_0372_);
  assign _0374_ = _0373_ ^ _0370_;
  assign _0375_ = b_i[12] & a_i[11];
  assign _0376_ = b_i[13] & a_i[10];
  assign _0377_ = ~(_0376_ ^ _0375_);
  assign _0378_ = b_i[14] & a_i[9];
  assign _0379_ = _0378_ ^ _0377_;
  assign _0380_ = _0379_ ^ _0374_;
  assign _0381_ = _0380_ ^ _0364_;
  assign _0382_ = _0308_ | _0305_;
  assign _0383_ = _0309_ & ~(_0315_);
  assign _0384_ = _0382_ & ~(_0383_);
  assign _0385_ = _0384_ ^ _0381_;
  assign _0386_ = _0385_ ^ _0363_;
  assign _0387_ = _0298_ & ~(_0321_);
  assign _0389_ = _0387_ ^ _0386_;
  assign _0390_ = ~_0389_;
  assign _0391_ = _0316_ | _0299_;
  assign _0392_ = _0317_ & ~(_0320_);
  assign _0393_ = _0391_ & ~(_0392_);
  assign _0394_ = ~(_0311_ & _0310_);
  assign _0395_ = _0314_ & ~(_0312_);
  assign _0396_ = _0394_ & ~(_0395_);
  assign _0397_ = ~(_0396_ ^ _0393_);
  assign _0398_ = b_i[15] & a_i[8];
  assign _0400_ = _0398_ ^ _0397_;
  assign _0401_ = _0400_ ^ _0390_;
  assign _0402_ = _0326_ | _0322_;
  assign _0403_ = ~(_0337_ | _0327_);
  assign _0404_ = _0402_ & ~(_0403_);
  assign _0405_ = ~(_0404_ ^ _0401_);
  assign _0406_ = _0333_ | _0330_;
  assign _0407_ = _0336_ & ~(_0334_);
  assign _0408_ = _0406_ & ~(_0407_);
  assign _0409_ = ~(_0408_ ^ _0405_);
  assign _0411_ = ~_0409_;
  assign _0412_ = _0341_ | _0338_;
  assign _0413_ = _0342_ & ~(_0345_);
  assign _0414_ = _0412_ & ~(_0413_);
  assign _0415_ = _0414_ ^ _0411_;
  assign _0416_ = _0350_ | _0347_;
  assign _0417_ = ~(_0358_ | _0351_);
  assign _0418_ = _0416_ & ~(_0417_);
  assign o[23] = _0418_ ^ _0415_;
  assign _0419_ = _0361_ & ~(_0360_);
  assign _0421_ = b_i[9] & a_i[15];
  assign _0422_ = b_i[10] & a_i[14];
  assign _0423_ = ~(_0422_ ^ _0421_);
  assign _0424_ = b_i[11] & a_i[13];
  assign _0425_ = _0424_ ^ _0423_;
  assign _0426_ = ~(_0366_ & _0365_);
  assign _0427_ = _0369_ & ~(_0368_);
  assign _0428_ = _0426_ & ~(_0427_);
  assign _0429_ = _0428_ ^ _0425_;
  assign _0430_ = b_i[12] & a_i[12];
  assign _0432_ = b_i[13] & a_i[11];
  assign _0433_ = ~(_0432_ ^ _0430_);
  assign _0434_ = b_i[14] & a_i[10];
  assign _0435_ = _0434_ ^ _0433_;
  assign _0436_ = _0435_ ^ _0429_;
  assign _0437_ = _0436_ ^ _0419_;
  assign _0438_ = _0373_ | _0370_;
  assign _0439_ = _0374_ & ~(_0379_);
  assign _0440_ = _0438_ & ~(_0439_);
  assign _0441_ = ~(_0440_ ^ _0437_);
  assign _0443_ = _0363_ & ~(_0385_);
  assign _0444_ = _0443_ ^ _0441_;
  assign _0445_ = ~_0444_;
  assign _0446_ = _0380_ | _0364_;
  assign _0447_ = _0381_ & ~(_0384_);
  assign _0448_ = _0446_ & ~(_0447_);
  assign _0449_ = ~(_0376_ & _0375_);
  assign _0450_ = _0378_ & ~(_0377_);
  assign _0451_ = _0449_ & ~(_0450_);
  assign _0452_ = ~(_0451_ ^ _0448_);
  assign _0454_ = b_i[15] & a_i[9];
  assign _0455_ = _0454_ ^ _0452_;
  assign _0456_ = _0455_ ^ _0445_;
  assign _0457_ = _0386_ | ~(_0387_);
  assign _0458_ = _0390_ & ~(_0400_);
  assign _0459_ = _0457_ & ~(_0458_);
  assign _0460_ = ~(_0459_ ^ _0456_);
  assign _0461_ = _0396_ | _0393_;
  assign _0462_ = _0398_ & ~(_0397_);
  assign _0463_ = _0461_ & ~(_0462_);
  assign _0465_ = ~(_0463_ ^ _0460_);
  assign _0466_ = _0404_ | _0401_;
  assign _0467_ = ~(_0408_ | _0405_);
  assign _0468_ = _0466_ & ~(_0467_);
  assign _0469_ = ~(_0468_ ^ _0465_);
  assign _0470_ = _0411_ & ~(_0414_);
  assign _0471_ = ~(_0416_ | _0415_);
  assign _0472_ = _0471_ | _0470_;
  assign _0473_ = _0415_ | _0351_;
  assign _0474_ = _0354_ & ~(_0473_);
  assign _0476_ = _0474_ | _0472_;
  assign _0477_ = _0473_ | _0355_;
  assign _0478_ = _0213_ & ~(_0477_);
  assign _0479_ = _0478_ | _0476_;
  assign _0480_ = _0477_ | _0214_;
  assign _0481_ = _1413_ & ~(_0480_);
  assign _0482_ = _0481_ | _0479_;
  assign o[24] = ~(_0482_ ^ _0469_);
  assign _0483_ = b_i[10] & a_i[15];
  assign _0484_ = b_i[11] & a_i[14];
  assign _0486_ = ~(_0484_ ^ _0483_);
  assign _0487_ = ~(_0422_ & _0421_);
  assign _0488_ = _0424_ & ~(_0423_);
  assign _0489_ = _0487_ & ~(_0488_);
  assign _0490_ = ~(_0489_ ^ _0486_);
  assign _0491_ = b_i[12] & a_i[13];
  assign _0492_ = b_i[13] & a_i[12];
  assign _0493_ = ~(_0492_ ^ _0491_);
  assign _0494_ = b_i[14] & a_i[11];
  assign _0495_ = _0494_ ^ _0493_;
  assign _0497_ = ~(_0495_ ^ _0490_);
  assign _0498_ = ~_0497_;
  assign _0499_ = _0428_ | _0425_;
  assign _0500_ = _0429_ & ~(_0435_);
  assign _0501_ = _0499_ & ~(_0500_);
  assign _0502_ = _0501_ ^ _0498_;
  assign _0503_ = ~_0502_;
  assign _0504_ = _0436_ | ~(_0419_);
  assign _0505_ = ~(_0440_ | _0437_);
  assign _0506_ = _0504_ & ~(_0505_);
  assign _0508_ = ~(_0432_ & _0430_);
  assign _0509_ = _0434_ & ~(_0433_);
  assign _0510_ = _0508_ & ~(_0509_);
  assign _0511_ = ~(_0510_ ^ _0506_);
  assign _0512_ = b_i[15] & a_i[10];
  assign _0513_ = _0512_ ^ _0511_;
  assign _0514_ = _0513_ ^ _0503_;
  assign _0515_ = _0441_ | ~(_0443_);
  assign _0516_ = _0445_ & ~(_0455_);
  assign _0517_ = _0515_ & ~(_0516_);
  assign _0519_ = ~(_0517_ ^ _0514_);
  assign _0520_ = _0451_ | _0448_;
  assign _0521_ = _0454_ & ~(_0452_);
  assign _0522_ = _0520_ & ~(_0521_);
  assign _0523_ = ~(_0522_ ^ _0519_);
  assign _0524_ = ~_0523_;
  assign _0525_ = _0459_ | _0456_;
  assign _0526_ = ~(_0463_ | _0460_);
  assign _0527_ = _0525_ & ~(_0526_);
  assign _0528_ = _0527_ ^ _0524_;
  assign _0530_ = _0468_ | _0465_;
  assign _0531_ = _0482_ & ~(_0469_);
  assign _0532_ = _0530_ & ~(_0531_);
  assign o[25] = _0532_ ^ _0528_;
  assign _0533_ = b_i[11] & a_i[15];
  assign _0534_ = _0484_ & _0483_;
  assign _0535_ = ~(_0534_ ^ _0533_);
  assign _0536_ = b_i[12] & a_i[14];
  assign _0537_ = b_i[13] & a_i[13];
  assign _0538_ = ~(_0537_ ^ _0536_);
  assign _0540_ = b_i[14] & a_i[12];
  assign _0541_ = _0540_ ^ _0538_;
  assign _0542_ = ~(_0541_ ^ _0535_);
  assign _0543_ = ~_0542_;
  assign _0544_ = _0489_ | _0486_;
  assign _0545_ = ~(_0495_ | _0490_);
  assign _0546_ = _0544_ & ~(_0545_);
  assign _0547_ = _0546_ ^ _0543_;
  assign _0548_ = ~_0547_;
  assign _0549_ = _0498_ & ~(_0501_);
  assign _0551_ = ~(_0492_ & _0491_);
  assign _0552_ = _0494_ & ~(_0493_);
  assign _0553_ = _0551_ & ~(_0552_);
  assign _0554_ = _0553_ ^ _0549_;
  assign _0555_ = b_i[15] & a_i[11];
  assign _0556_ = _0555_ ^ _0554_;
  assign _0557_ = _0556_ ^ _0548_;
  assign _0558_ = _0503_ & ~(_0513_);
  assign _0559_ = _0558_ ^ _0557_;
  assign _0560_ = _0510_ | _0506_;
  assign _0562_ = _0512_ & ~(_0511_);
  assign _0563_ = _0560_ & ~(_0562_);
  assign _0564_ = ~(_0563_ ^ _0559_);
  assign _0565_ = _0517_ | _0514_;
  assign _0566_ = ~(_0522_ | _0519_);
  assign _0567_ = _0565_ & ~(_0566_);
  assign _0568_ = ~(_0567_ ^ _0564_);
  assign _0569_ = _0524_ & ~(_0527_);
  assign _0570_ = ~(_0530_ | _0528_);
  assign _0571_ = ~(_0570_ | _0569_);
  assign _0573_ = _0528_ | _0469_;
  assign _0574_ = _0482_ & ~(_0573_);
  assign _0575_ = _0571_ & ~(_0574_);
  assign o[26] = _0575_ ^ _0568_;
  assign _0576_ = b_i[12] & a_i[15];
  assign _0577_ = b_i[13] & a_i[14];
  assign _0578_ = ~(_0577_ ^ _0576_);
  assign _0579_ = b_i[14] & a_i[13];
  assign _0580_ = _0579_ ^ _0578_;
  assign _0581_ = ~_0580_;
  assign _0583_ = ~(_0534_ & _0533_);
  assign _0584_ = ~(_0541_ | _0535_);
  assign _0585_ = _0583_ & ~(_0584_);
  assign _0586_ = _0585_ ^ _0581_;
  assign _0587_ = ~_0586_;
  assign _0588_ = _0543_ & ~(_0546_);
  assign _0589_ = ~(_0537_ & _0536_);
  assign _0590_ = _0540_ & ~(_0538_);
  assign _0591_ = _0589_ & ~(_0590_);
  assign _0592_ = _0591_ ^ _0588_;
  assign _0594_ = b_i[15] & a_i[12];
  assign _0595_ = _0594_ ^ _0592_;
  assign _0596_ = _0595_ ^ _0587_;
  assign _0597_ = _0548_ & ~(_0556_);
  assign _0598_ = _0597_ ^ _0596_;
  assign _0599_ = _0553_ | ~(_0549_);
  assign _0600_ = _0555_ & ~(_0554_);
  assign _0601_ = _0599_ & ~(_0600_);
  assign _0602_ = ~(_0601_ ^ _0598_);
  assign _0603_ = _0557_ | ~(_0558_);
  assign _0605_ = ~(_0563_ | _0559_);
  assign _0606_ = _0603_ & ~(_0605_);
  assign _0607_ = ~(_0606_ ^ _0602_);
  assign _0608_ = _0567_ | _0564_;
  assign _0609_ = ~(_0575_ | _0568_);
  assign _0610_ = _0608_ & ~(_0609_);
  assign o[27] = _0610_ ^ _0607_;
  assign _0611_ = b_i[13] & a_i[15];
  assign _0612_ = b_i[14] & a_i[14];
  assign _0613_ = ~(_0612_ ^ _0611_);
  assign _0615_ = ~_0613_;
  assign _0616_ = _0581_ & ~(_0585_);
  assign _0617_ = ~(_0577_ & _0576_);
  assign _0618_ = _0579_ & ~(_0578_);
  assign _0619_ = _0617_ & ~(_0618_);
  assign _0620_ = _0619_ ^ _0616_;
  assign _0621_ = b_i[15] & a_i[13];
  assign _0622_ = _0621_ ^ _0620_;
  assign _0623_ = _0622_ ^ _0615_;
  assign _0624_ = _0587_ & ~(_0595_);
  assign _0626_ = _0624_ ^ _0623_;
  assign _0627_ = _0591_ | ~(_0588_);
  assign _0628_ = _0594_ & ~(_0592_);
  assign _0629_ = _0627_ & ~(_0628_);
  assign _0630_ = ~(_0629_ ^ _0626_);
  assign _0631_ = _0596_ | ~(_0597_);
  assign _0632_ = ~(_0601_ | _0598_);
  assign _0633_ = _0631_ & ~(_0632_);
  assign _0634_ = ~(_0633_ ^ _0630_);
  assign _0635_ = _0606_ | _0602_;
  assign _0637_ = ~(_0608_ | _0607_);
  assign _0638_ = _0635_ & ~(_0637_);
  assign _0639_ = _0607_ | _0568_;
  assign _0640_ = ~(_0639_ | _0571_);
  assign _0641_ = _0638_ & ~(_0640_);
  assign _0642_ = _0639_ | _0573_;
  assign _0643_ = _0482_ & ~(_0642_);
  assign _0644_ = _0641_ & ~(_0643_);
  assign o[28] = _0644_ ^ _0634_;
  assign _0645_ = b_i[14] & a_i[15];
  assign _0647_ = _0612_ & _0611_;
  assign _0648_ = b_i[15] & a_i[14];
  assign _0649_ = ~_0648_;
  assign _0650_ = _0649_ ^ _0647_;
  assign _0651_ = _0650_ ^ _0645_;
  assign _0652_ = _0615_ & ~(_0622_);
  assign _0653_ = _0652_ ^ _0651_;
  assign _0654_ = _0619_ | ~(_0616_);
  assign _0655_ = _0621_ & ~(_0620_);
  assign _0656_ = _0654_ & ~(_0655_);
  assign _0658_ = ~(_0656_ ^ _0653_);
  assign _0659_ = _0623_ | ~(_0624_);
  assign _0660_ = ~(_0629_ | _0626_);
  assign _0661_ = _0659_ & ~(_0660_);
  assign _0662_ = ~(_0661_ ^ _0658_);
  assign _0663_ = _0633_ | _0630_;
  assign _0664_ = ~(_0644_ | _0634_);
  assign _0665_ = _0663_ & ~(_0664_);
  assign o[29] = _0665_ ^ _0662_;
  assign _0666_ = b_i[15] & a_i[15];
  assign _0668_ = _0645_ & ~(_0650_);
  assign _0669_ = ~(_0668_ ^ _0666_);
  assign _0670_ = _0647_ & ~(_0649_);
  assign _0671_ = _0670_ ^ _0669_;
  assign _0672_ = _0651_ | ~(_0652_);
  assign _0673_ = ~(_0656_ | _0653_);
  assign _0674_ = _0672_ & ~(_0673_);
  assign _0675_ = ~(_0674_ ^ _0671_);
  assign _0676_ = _0661_ | _0658_;
  assign _0677_ = ~(_0663_ | _0662_);
  assign _0679_ = _0676_ & ~(_0677_);
  assign _0680_ = _0662_ | _0634_;
  assign _0681_ = ~(_0680_ | _0644_);
  assign _0682_ = _0679_ & ~(_0681_);
  assign o[30] = _0682_ ^ _0675_;
  assign _0683_ = ~(_0668_ & _0666_);
  assign _0684_ = _0670_ & ~(_0669_);
  assign _0685_ = _0683_ & ~(_0684_);
  assign _0686_ = _0674_ | _0671_;
  assign _0687_ = ~(_0682_ | _0675_);
  assign _0689_ = _0686_ & ~(_0687_);
  assign o[31] = _0689_ ^ _0685_;
  assign o[7] = ~(_0780_ ^ _0779_);
  assign o[1] = _1254_ ^ _1243_;
endmodule
