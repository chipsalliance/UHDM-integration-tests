module bsg_decode(i, o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  input [3:0] i;
  wire [3:0] i;
  output [15:0] o;
  wire [15:0] o;
  assign _00_ = ~i[3];
  assign _01_ = i[0] | i[1];
  assign _02_ = _01_ | i[2];
  assign o[0] = _00_ & ~(_02_);
  assign _03_ = i[1] | ~(i[0]);
  assign _04_ = _03_ | i[2];
  assign o[1] = _00_ & ~(_04_);
  assign _05_ = i[0] | ~(i[1]);
  assign _06_ = _05_ | i[2];
  assign o[2] = _00_ & ~(_06_);
  assign _07_ = ~(i[0] & i[1]);
  assign _08_ = _07_ | i[2];
  assign o[3] = _00_ & ~(_08_);
  assign _09_ = ~i[2];
  assign _10_ = _01_ | _09_;
  assign o[4] = _00_ & ~(_10_);
  assign _11_ = _03_ | _09_;
  assign o[5] = _00_ & ~(_11_);
  assign _12_ = _05_ | _09_;
  assign o[6] = _00_ & ~(_12_);
  assign _13_ = _07_ | _09_;
  assign o[7] = _00_ & ~(_13_);
  assign o[8] = i[3] & ~(_02_);
  assign o[9] = i[3] & ~(_04_);
  assign o[10] = i[3] & ~(_06_);
  assign o[11] = i[3] & ~(_08_);
  assign o[12] = i[3] & ~(_10_);
  assign o[13] = i[3] & ~(_11_);
  assign o[14] = i[3] & ~(_12_);
  assign o[15] = i[3] & ~(_13_);
endmodule
