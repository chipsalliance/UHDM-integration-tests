module bsg_fsb_node_async_buffer(L_clk_i, L_reset_i, L_en_o, L_v_o, L_data_o, L_ready_i, L_v_i, L_data_i, L_yumi_o, R_clk_i, R_reset_i, R_en_i, R_v_i, R_data_i, R_ready_o, R_v_o, R_data_o, R_yumi_i);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  input L_clk_i;
  wire L_clk_i;
  input [4:0] L_data_i;
  wire [4:0] L_data_i;
  output [4:0] L_data_o;
  wire [4:0] L_data_o;
  output L_en_o;
  wire L_en_o;
  input L_ready_i;
  wire L_ready_i;
  input L_reset_i;
  wire L_reset_i;
  input L_v_i;
  wire L_v_i;
  output L_v_o;
  wire L_v_o;
  wire L_w_full_lo;
  output L_yumi_o;
  wire L_yumi_o;
  input R_clk_i;
  wire R_clk_i;
  input [4:0] R_data_i;
  wire [4:0] R_data_i;
  output [4:0] R_data_o;
  wire [4:0] R_data_o;
  input R_en_i;
  wire R_en_i;
  output R_ready_o;
  wire R_ready_o;
  input R_reset_i;
  wire R_reset_i;
  input R_v_i;
  wire R_v_i;
  output R_v_o;
  wire R_v_o;
  wire R_w_full_lo;
  input R_yumi_i;
  wire R_yumi_i;
  wire \fsb_en_sync.iclk_data_i ;
  wire \fsb_en_sync.oclk_data_o ;
  wire \fsb_en_sync.oclk_i ;
  reg \fsb_en_sync.z.bss.bsg_SYNC_1_r ;
  reg \fsb_en_sync.z.bss.bsg_SYNC_2_r ;
  wire \fsb_en_sync.z.bss.iclk_data_i ;
  wire \fsb_en_sync.z.bss.oclk_data_o ;
  wire \fsb_en_sync.z.bss.oclk_i ;
  wire \l2r_fifo.MSYNC_1r1w.r_addr_i ;
  wire [4:0] \l2r_fifo.MSYNC_1r1w.r_data_o ;
  wire \l2r_fifo.MSYNC_1r1w.r_v_i ;
  reg [4:0] \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] ;
  reg [4:0] \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] ;
  wire \l2r_fifo.MSYNC_1r1w.synth.r_addr_i ;
  wire [4:0] \l2r_fifo.MSYNC_1r1w.synth.r_data_o ;
  wire \l2r_fifo.MSYNC_1r1w.synth.r_v_i ;
  wire \l2r_fifo.MSYNC_1r1w.synth.unused0 ;
  wire \l2r_fifo.MSYNC_1r1w.synth.unused1 ;
  wire \l2r_fifo.MSYNC_1r1w.synth.w_addr_i ;
  wire \l2r_fifo.MSYNC_1r1w.synth.w_clk_i ;
  wire [4:0] \l2r_fifo.MSYNC_1r1w.synth.w_data_i ;
  wire \l2r_fifo.MSYNC_1r1w.synth.w_reset_i ;
  wire \l2r_fifo.MSYNC_1r1w.synth.w_v_i ;
  wire \l2r_fifo.MSYNC_1r1w.w_addr_i ;
  wire \l2r_fifo.MSYNC_1r1w.w_clk_i ;
  wire [4:0] \l2r_fifo.MSYNC_1r1w.w_data_i ;
  wire \l2r_fifo.MSYNC_1r1w.w_reset_i ;
  wire \l2r_fifo.MSYNC_1r1w.w_v_i ;
  wire [1:0] \l2r_fifo.bapg_rd.ptr_sync.iclk_data_o ;
  wire \l2r_fifo.bapg_rd.ptr_sync.iclk_i ;
  wire \l2r_fifo.bapg_rd.ptr_sync.iclk_reset_i ;
  wire [1:0] \l2r_fifo.bapg_rd.ptr_sync.oclk_data_o ;
  wire \l2r_fifo.bapg_rd.ptr_sync.oclk_i ;
  reg [1:0] \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r ;
  reg [1:0] \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  reg [1:0] \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  wire [1:0] \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_data_o ;
  wire \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_i ;
  wire \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_reset_i ;
  wire [1:0] \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.oclk_data_o ;
  wire \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.oclk_i ;
  wire \l2r_fifo.bapg_rd.r_clk_i ;
  wire \l2r_fifo.bapg_rd.w_clk_i ;
  wire \l2r_fifo.bapg_rd.w_inc_i ;
  wire [1:0] \l2r_fifo.bapg_rd.w_ptr_binary_r_o ;
  wire [1:0] \l2r_fifo.bapg_rd.w_ptr_gray_r ;
  wire [1:0] \l2r_fifo.bapg_rd.w_ptr_gray_r_o ;
  wire [1:0] \l2r_fifo.bapg_rd.w_ptr_gray_r_rsync ;
  wire [1:0] \l2r_fifo.bapg_rd.w_ptr_gray_r_rsync_o ;
  wire [1:0] \l2r_fifo.bapg_rd.w_ptr_p1_r ;
  wire [1:0] \l2r_fifo.bapg_rd.w_ptr_p2 ;
  wire [1:0] \l2r_fifo.bapg_rd.w_ptr_r ;
  wire \l2r_fifo.bapg_rd.w_reset_i ;
  wire [1:0] \l2r_fifo.bapg_wr.ptr_sync.iclk_data_o ;
  wire \l2r_fifo.bapg_wr.ptr_sync.iclk_i ;
  wire \l2r_fifo.bapg_wr.ptr_sync.iclk_reset_i ;
  wire [1:0] \l2r_fifo.bapg_wr.ptr_sync.oclk_data_o ;
  wire \l2r_fifo.bapg_wr.ptr_sync.oclk_i ;
  reg [1:0] \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r ;
  reg [1:0] \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  reg [1:0] \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  wire [1:0] \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_data_o ;
  wire \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_i ;
  wire \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_reset_i ;
  wire [1:0] \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.oclk_data_o ;
  wire \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.oclk_i ;
  wire \l2r_fifo.bapg_wr.r_clk_i ;
  wire \l2r_fifo.bapg_wr.w_clk_i ;
  wire \l2r_fifo.bapg_wr.w_inc_i ;
  wire [1:0] \l2r_fifo.bapg_wr.w_ptr_binary_r_o ;
  wire [1:0] \l2r_fifo.bapg_wr.w_ptr_gray_r ;
  wire [1:0] \l2r_fifo.bapg_wr.w_ptr_gray_r_o ;
  wire [1:0] \l2r_fifo.bapg_wr.w_ptr_gray_r_rsync ;
  wire [1:0] \l2r_fifo.bapg_wr.w_ptr_gray_r_rsync_o ;
  wire [1:0] \l2r_fifo.bapg_wr.w_ptr_p1_r ;
  wire [1:0] \l2r_fifo.bapg_wr.w_ptr_p2 ;
  wire [1:0] \l2r_fifo.bapg_wr.w_ptr_r ;
  wire \l2r_fifo.bapg_wr.w_reset_i ;
  wire \l2r_fifo.r_clk_i ;
  wire [4:0] \l2r_fifo.r_data_o ;
  wire [4:0] \l2r_fifo.r_data_o_tmp ;
  wire \l2r_fifo.r_deq_i ;
  wire [1:0] \l2r_fifo.r_ptr_binary_r ;
  wire [1:0] \l2r_fifo.r_ptr_gray_r ;
  wire [1:0] \l2r_fifo.r_ptr_gray_r_wsync ;
  wire \l2r_fifo.r_reset_i ;
  wire \l2r_fifo.r_valid_o ;
  wire \l2r_fifo.r_valid_o_tmp ;
  wire \l2r_fifo.w_clk_i ;
  wire [4:0] \l2r_fifo.w_data_i ;
  wire \l2r_fifo.w_enq_i ;
  wire \l2r_fifo.w_full_o ;
  wire [1:0] \l2r_fifo.w_ptr_binary_r ;
  wire [1:0] \l2r_fifo.w_ptr_gray_r ;
  wire [1:0] \l2r_fifo.w_ptr_gray_r_rsync ;
  wire \l2r_fifo.w_reset_i ;
  wire \r2l_fifo.MSYNC_1r1w.r_addr_i ;
  wire [4:0] \r2l_fifo.MSYNC_1r1w.r_data_o ;
  wire \r2l_fifo.MSYNC_1r1w.r_v_i ;
  reg [4:0] \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] ;
  reg [4:0] \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] ;
  wire \r2l_fifo.MSYNC_1r1w.synth.r_addr_i ;
  wire [4:0] \r2l_fifo.MSYNC_1r1w.synth.r_data_o ;
  wire \r2l_fifo.MSYNC_1r1w.synth.r_v_i ;
  wire \r2l_fifo.MSYNC_1r1w.synth.unused0 ;
  wire \r2l_fifo.MSYNC_1r1w.synth.unused1 ;
  wire \r2l_fifo.MSYNC_1r1w.synth.w_addr_i ;
  wire \r2l_fifo.MSYNC_1r1w.synth.w_clk_i ;
  wire [4:0] \r2l_fifo.MSYNC_1r1w.synth.w_data_i ;
  wire \r2l_fifo.MSYNC_1r1w.synth.w_reset_i ;
  wire \r2l_fifo.MSYNC_1r1w.synth.w_v_i ;
  wire \r2l_fifo.MSYNC_1r1w.w_addr_i ;
  wire \r2l_fifo.MSYNC_1r1w.w_clk_i ;
  wire [4:0] \r2l_fifo.MSYNC_1r1w.w_data_i ;
  wire \r2l_fifo.MSYNC_1r1w.w_reset_i ;
  wire \r2l_fifo.MSYNC_1r1w.w_v_i ;
  wire [1:0] \r2l_fifo.bapg_rd.ptr_sync.iclk_data_o ;
  wire \r2l_fifo.bapg_rd.ptr_sync.iclk_i ;
  wire \r2l_fifo.bapg_rd.ptr_sync.iclk_reset_i ;
  wire [1:0] \r2l_fifo.bapg_rd.ptr_sync.oclk_data_o ;
  wire \r2l_fifo.bapg_rd.ptr_sync.oclk_i ;
  reg [1:0] \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r ;
  reg [1:0] \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  reg [1:0] \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  wire [1:0] \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_data_o ;
  wire \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_i ;
  wire \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_reset_i ;
  wire [1:0] \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.oclk_data_o ;
  wire \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.oclk_i ;
  wire \r2l_fifo.bapg_rd.r_clk_i ;
  wire \r2l_fifo.bapg_rd.w_clk_i ;
  wire \r2l_fifo.bapg_rd.w_inc_i ;
  wire [1:0] \r2l_fifo.bapg_rd.w_ptr_binary_r_o ;
  wire [1:0] \r2l_fifo.bapg_rd.w_ptr_gray_r ;
  wire [1:0] \r2l_fifo.bapg_rd.w_ptr_gray_r_o ;
  wire [1:0] \r2l_fifo.bapg_rd.w_ptr_gray_r_rsync ;
  wire [1:0] \r2l_fifo.bapg_rd.w_ptr_gray_r_rsync_o ;
  wire [1:0] \r2l_fifo.bapg_rd.w_ptr_p1_r ;
  wire [1:0] \r2l_fifo.bapg_rd.w_ptr_p2 ;
  wire [1:0] \r2l_fifo.bapg_rd.w_ptr_r ;
  wire \r2l_fifo.bapg_rd.w_reset_i ;
  wire [1:0] \r2l_fifo.bapg_wr.ptr_sync.iclk_data_o ;
  wire \r2l_fifo.bapg_wr.ptr_sync.iclk_i ;
  wire \r2l_fifo.bapg_wr.ptr_sync.iclk_reset_i ;
  wire [1:0] \r2l_fifo.bapg_wr.ptr_sync.oclk_data_o ;
  wire \r2l_fifo.bapg_wr.ptr_sync.oclk_i ;
  reg [1:0] \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r ;
  reg [1:0] \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  reg [1:0] \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  wire [1:0] \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_data_o ;
  wire \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_i ;
  wire \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_reset_i ;
  wire [1:0] \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.oclk_data_o ;
  wire \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.oclk_i ;
  wire \r2l_fifo.bapg_wr.r_clk_i ;
  wire \r2l_fifo.bapg_wr.w_clk_i ;
  wire \r2l_fifo.bapg_wr.w_inc_i ;
  wire [1:0] \r2l_fifo.bapg_wr.w_ptr_binary_r_o ;
  wire [1:0] \r2l_fifo.bapg_wr.w_ptr_gray_r ;
  wire [1:0] \r2l_fifo.bapg_wr.w_ptr_gray_r_o ;
  wire [1:0] \r2l_fifo.bapg_wr.w_ptr_gray_r_rsync ;
  wire [1:0] \r2l_fifo.bapg_wr.w_ptr_gray_r_rsync_o ;
  wire [1:0] \r2l_fifo.bapg_wr.w_ptr_p1_r ;
  wire [1:0] \r2l_fifo.bapg_wr.w_ptr_p2 ;
  wire [1:0] \r2l_fifo.bapg_wr.w_ptr_r ;
  wire \r2l_fifo.bapg_wr.w_reset_i ;
  wire \r2l_fifo.r_clk_i ;
  wire [4:0] \r2l_fifo.r_data_o ;
  wire [4:0] \r2l_fifo.r_data_o_tmp ;
  wire \r2l_fifo.r_deq_i ;
  wire [1:0] \r2l_fifo.r_ptr_binary_r ;
  wire [1:0] \r2l_fifo.r_ptr_gray_r ;
  wire [1:0] \r2l_fifo.r_ptr_gray_r_wsync ;
  wire \r2l_fifo.r_reset_i ;
  wire \r2l_fifo.r_valid_o ;
  wire \r2l_fifo.r_valid_o_tmp ;
  wire \r2l_fifo.w_clk_i ;
  wire [4:0] \r2l_fifo.w_data_i ;
  wire \r2l_fifo.w_enq_i ;
  wire \r2l_fifo.w_full_o ;
  wire [1:0] \r2l_fifo.w_ptr_binary_r ;
  wire [1:0] \r2l_fifo.w_ptr_gray_r ;
  wire [1:0] \r2l_fifo.w_ptr_gray_r_rsync ;
  wire \r2l_fifo.w_reset_i ;
  assign \l2r_fifo.bapg_rd.w_ptr_p2 [0] = ~\l2r_fifo.bapg_rd.w_ptr_p1_r [0];
  assign \r2l_fifo.bapg_wr.w_ptr_p2 [0] = ~\r2l_fifo.bapg_wr.w_ptr_p1_r [0];
  assign _007_ = ~(\r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] ^ \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0]);
  assign _008_ = ~(\r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] & \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0]);
  assign R_ready_o = _008_ | ~(_007_);
  assign _009_ = ~(\r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] ^ \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0]);
  assign _010_ = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] ^ \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1];
  assign L_v_o = _010_ | ~(_009_);
  assign _011_ = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] ^ \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  assign _012_ = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] ^ \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1];
  assign R_v_o = _012_ | _011_;
  assign L_data_o[0] = \r2l_fifo.bapg_rd.w_ptr_r [0] ? \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [0] : \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [0];
  assign L_data_o[1] = \r2l_fifo.bapg_rd.w_ptr_r [0] ? \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [1] : \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [1];
  assign L_data_o[2] = \r2l_fifo.bapg_rd.w_ptr_r [0] ? \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [2] : \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [2];
  assign L_data_o[3] = \r2l_fifo.bapg_rd.w_ptr_r [0] ? \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [3] : \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [3];
  assign L_data_o[4] = \r2l_fifo.bapg_rd.w_ptr_r [0] ? \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [4] : \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [4];
  assign R_data_o[0] = \l2r_fifo.bapg_rd.w_ptr_r [0] ? \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [0] : \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [0];
  assign R_data_o[1] = \l2r_fifo.bapg_rd.w_ptr_r [0] ? \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [1] : \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [1];
  assign R_data_o[2] = \l2r_fifo.bapg_rd.w_ptr_r [0] ? \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [2] : \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [2];
  assign R_data_o[3] = \l2r_fifo.bapg_rd.w_ptr_r [0] ? \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [3] : \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [3];
  assign R_data_o[4] = \l2r_fifo.bapg_rd.w_ptr_r [0] ? \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [4] : \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [4];
  assign \r2l_fifo.bapg_rd.w_ptr_p2 [0] = ~\r2l_fifo.bapg_rd.w_ptr_p1_r [0];
  assign \l2r_fifo.bapg_wr.w_ptr_p2 [0] = ~\l2r_fifo.bapg_wr.w_ptr_p1_r [0];
  assign \r2l_fifo.bapg_wr.w_inc_i  = R_ready_o & R_v_i;
  assign \r2l_fifo.bapg_rd.w_inc_i  = L_v_o & L_ready_i;
  assign _004_ = ~(\l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] ^ \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0]);
  assign _005_ = ~(\l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] & \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0]);
  assign _006_ = _004_ & ~(_005_);
  assign \l2r_fifo.bapg_wr.w_inc_i  = L_v_i & ~(_006_);
  assign _003_ = \r2l_fifo.bapg_wr.w_inc_i  & \r2l_fifo.bapg_wr.w_ptr_r [0];
  assign _000_ = \l2r_fifo.bapg_wr.w_inc_i  & ~(\l2r_fifo.bapg_wr.w_ptr_r [0]);
  assign _002_ = \r2l_fifo.bapg_wr.w_inc_i  & ~(\r2l_fifo.bapg_wr.w_ptr_r [0]);
  assign _001_ = \l2r_fifo.bapg_wr.w_inc_i  & \l2r_fifo.bapg_wr.w_ptr_r [0];
  assign \l2r_fifo.bapg_rd.w_ptr_p2 [1] = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] ^ \l2r_fifo.bapg_rd.w_ptr_p1_r [0];
  assign \r2l_fifo.bapg_rd.w_ptr_p2 [1] = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] ^ \r2l_fifo.bapg_rd.w_ptr_p1_r [0];
  assign \r2l_fifo.bapg_wr.w_ptr_p2 [1] = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] ^ \r2l_fifo.bapg_wr.w_ptr_p1_r [0];
  assign \l2r_fifo.bapg_wr.w_ptr_p2 [1] = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] ^ \l2r_fifo.bapg_wr.w_ptr_p1_r [0];
  always @(posedge R_clk_i)
    if (_002_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [0] <= R_data_i[0];
  always @(posedge R_clk_i)
    if (_002_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [1] <= R_data_i[1];
  always @(posedge R_clk_i)
    if (_002_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [2] <= R_data_i[2];
  always @(posedge R_clk_i)
    if (_002_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [3] <= R_data_i[3];
  always @(posedge R_clk_i)
    if (_002_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[0] [4] <= R_data_i[4];
  always @(posedge R_clk_i)
    if (_003_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [0] <= R_data_i[0];
  always @(posedge R_clk_i)
    if (_003_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [1] <= R_data_i[1];
  always @(posedge R_clk_i)
    if (_003_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [2] <= R_data_i[2];
  always @(posedge R_clk_i)
    if (_003_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [3] <= R_data_i[3];
  always @(posedge R_clk_i)
    if (_003_) \r2l_fifo.MSYNC_1r1w.synth.nz.mem[1] [4] <= R_data_i[4];
  reg \r2l_fifo.bapg_rd.w_ptr_p1_r_reg[0] ;
  always @(posedge L_clk_i)
    if (L_reset_i) \r2l_fifo.bapg_rd.w_ptr_p1_r_reg[0]  <= 1'h1;
    else if (\r2l_fifo.bapg_rd.w_inc_i ) \r2l_fifo.bapg_rd.w_ptr_p1_r_reg[0]  <= \r2l_fifo.bapg_rd.w_ptr_p2 [0];
  assign \r2l_fifo.bapg_rd.w_ptr_p1_r [0] = \r2l_fifo.bapg_rd.w_ptr_p1_r_reg[0] ;
  reg \r2l_fifo.bapg_rd.w_ptr_r_reg[0] ;
  always @(posedge L_clk_i)
    if (L_reset_i) \r2l_fifo.bapg_rd.w_ptr_r_reg[0]  <= 1'h0;
    else if (\r2l_fifo.bapg_rd.w_inc_i ) \r2l_fifo.bapg_rd.w_ptr_r_reg[0]  <= \r2l_fifo.bapg_rd.w_ptr_p1_r [0];
  assign \r2l_fifo.bapg_rd.w_ptr_r [0] = \r2l_fifo.bapg_rd.w_ptr_r_reg[0] ;
  always @(posedge R_clk_i)
    \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] <= \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0];
  always @(posedge R_clk_i)
    \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] <= \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1];
  always @(posedge R_clk_i)
    \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0] <= \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  always @(posedge R_clk_i)
    \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1] <= \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1];
  always @(posedge L_clk_i)
    if (L_reset_i) \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= 1'h0;
    else if (\r2l_fifo.bapg_rd.w_inc_i ) \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= \r2l_fifo.bapg_rd.w_ptr_p2 [1];
  always @(posedge L_clk_i)
    if (L_reset_i) \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= 1'h0;
    else if (\r2l_fifo.bapg_rd.w_inc_i ) \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  reg \r2l_fifo.bapg_wr.w_ptr_p1_r_reg[0] ;
  always @(posedge R_clk_i)
    if (R_reset_i) \r2l_fifo.bapg_wr.w_ptr_p1_r_reg[0]  <= 1'h1;
    else if (\r2l_fifo.bapg_wr.w_inc_i ) \r2l_fifo.bapg_wr.w_ptr_p1_r_reg[0]  <= \r2l_fifo.bapg_wr.w_ptr_p2 [0];
  assign \r2l_fifo.bapg_wr.w_ptr_p1_r [0] = \r2l_fifo.bapg_wr.w_ptr_p1_r_reg[0] ;
  reg \r2l_fifo.bapg_wr.w_ptr_r_reg[0] ;
  always @(posedge R_clk_i)
    if (R_reset_i) \r2l_fifo.bapg_wr.w_ptr_r_reg[0]  <= 1'h0;
    else if (\r2l_fifo.bapg_wr.w_inc_i ) \r2l_fifo.bapg_wr.w_ptr_r_reg[0]  <= \r2l_fifo.bapg_wr.w_ptr_p1_r [0];
  assign \r2l_fifo.bapg_wr.w_ptr_r [0] = \r2l_fifo.bapg_wr.w_ptr_r_reg[0] ;
  always @(posedge L_clk_i)
    \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] <= \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0];
  always @(posedge L_clk_i)
    \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] <= \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1];
  always @(posedge L_clk_i)
    \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0] <= \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  always @(posedge L_clk_i)
    \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1] <= \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1];
  always @(posedge R_clk_i)
    if (R_reset_i) \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= 1'h0;
    else if (\r2l_fifo.bapg_wr.w_inc_i ) \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= \r2l_fifo.bapg_wr.w_ptr_p2 [1];
  always @(posedge R_clk_i)
    if (R_reset_i) \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= 1'h0;
    else if (\r2l_fifo.bapg_wr.w_inc_i ) \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  always @(posedge L_clk_i)
    if (_001_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [0] <= L_data_i[0];
  always @(posedge L_clk_i)
    if (_001_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [1] <= L_data_i[1];
  always @(posedge L_clk_i)
    if (_001_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [2] <= L_data_i[2];
  always @(posedge L_clk_i)
    if (_001_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [3] <= L_data_i[3];
  always @(posedge L_clk_i)
    if (_001_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[1] [4] <= L_data_i[4];
  reg \l2r_fifo.bapg_rd.w_ptr_p1_r_reg[0] ;
  always @(posedge R_clk_i)
    if (R_reset_i) \l2r_fifo.bapg_rd.w_ptr_p1_r_reg[0]  <= 1'h1;
    else if (R_yumi_i) \l2r_fifo.bapg_rd.w_ptr_p1_r_reg[0]  <= \l2r_fifo.bapg_rd.w_ptr_p2 [0];
  assign \l2r_fifo.bapg_rd.w_ptr_p1_r [0] = \l2r_fifo.bapg_rd.w_ptr_p1_r_reg[0] ;
  reg \l2r_fifo.bapg_rd.w_ptr_r_reg[0] ;
  always @(posedge R_clk_i)
    if (R_reset_i) \l2r_fifo.bapg_rd.w_ptr_r_reg[0]  <= 1'h0;
    else if (R_yumi_i) \l2r_fifo.bapg_rd.w_ptr_r_reg[0]  <= \l2r_fifo.bapg_rd.w_ptr_p1_r [0];
  assign \l2r_fifo.bapg_rd.w_ptr_r [0] = \l2r_fifo.bapg_rd.w_ptr_r_reg[0] ;
  always @(posedge L_clk_i)
    \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] <= \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0];
  always @(posedge L_clk_i)
    \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] <= \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1];
  always @(posedge L_clk_i)
    \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0] <= \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  always @(posedge L_clk_i)
    \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1] <= \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1];
  always @(posedge R_clk_i)
    if (R_reset_i) \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= 1'h0;
    else if (R_yumi_i) \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= \l2r_fifo.bapg_rd.w_ptr_p2 [1];
  always @(posedge R_clk_i)
    if (R_reset_i) \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= 1'h0;
    else if (R_yumi_i) \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  reg \l2r_fifo.bapg_wr.w_ptr_p1_r_reg[0] ;
  always @(posedge L_clk_i)
    if (L_reset_i) \l2r_fifo.bapg_wr.w_ptr_p1_r_reg[0]  <= 1'h1;
    else if (\l2r_fifo.bapg_wr.w_inc_i ) \l2r_fifo.bapg_wr.w_ptr_p1_r_reg[0]  <= \l2r_fifo.bapg_wr.w_ptr_p2 [0];
  assign \l2r_fifo.bapg_wr.w_ptr_p1_r [0] = \l2r_fifo.bapg_wr.w_ptr_p1_r_reg[0] ;
  reg \l2r_fifo.bapg_wr.w_ptr_r_reg[0] ;
  always @(posedge L_clk_i)
    if (L_reset_i) \l2r_fifo.bapg_wr.w_ptr_r_reg[0]  <= 1'h0;
    else if (\l2r_fifo.bapg_wr.w_inc_i ) \l2r_fifo.bapg_wr.w_ptr_r_reg[0]  <= \l2r_fifo.bapg_wr.w_ptr_p1_r [0];
  assign \l2r_fifo.bapg_wr.w_ptr_r [0] = \l2r_fifo.bapg_wr.w_ptr_r_reg[0] ;
  always @(posedge R_clk_i)
    \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] <= \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0];
  always @(posedge R_clk_i)
    \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] <= \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1];
  always @(posedge R_clk_i)
    \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0] <= \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  always @(posedge R_clk_i)
    \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1] <= \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1];
  always @(posedge L_clk_i)
    if (L_reset_i) \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= 1'h0;
    else if (\l2r_fifo.bapg_wr.w_inc_i ) \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= \l2r_fifo.bapg_wr.w_ptr_p2 [1];
  always @(posedge L_clk_i)
    if (L_reset_i) \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= 1'h0;
    else if (\l2r_fifo.bapg_wr.w_inc_i ) \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  always @(posedge L_clk_i)
    if (_000_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [0] <= L_data_i[0];
  always @(posedge L_clk_i)
    if (_000_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [1] <= L_data_i[1];
  always @(posedge L_clk_i)
    if (_000_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [2] <= L_data_i[2];
  always @(posedge L_clk_i)
    if (_000_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [3] <= L_data_i[3];
  always @(posedge L_clk_i)
    if (_000_) \l2r_fifo.MSYNC_1r1w.synth.nz.mem[0] [4] <= L_data_i[4];
  always @(posedge L_clk_i)
    \fsb_en_sync.z.bss.bsg_SYNC_1_r  <= R_en_i;
  always @(posedge L_clk_i)
    \fsb_en_sync.z.bss.bsg_SYNC_2_r  <= \fsb_en_sync.z.bss.bsg_SYNC_1_r ;
  assign L_en_o = \fsb_en_sync.z.bss.bsg_SYNC_2_r ;
  assign L_w_full_lo = \l2r_fifo.w_full_o ;
  assign L_yumi_o = \l2r_fifo.bapg_wr.w_inc_i ;
  assign R_w_full_lo = \r2l_fifo.w_full_o ;
  assign \fsb_en_sync.iclk_data_i  = R_en_i;
  assign \fsb_en_sync.oclk_data_o  = \fsb_en_sync.z.bss.bsg_SYNC_2_r ;
  assign \fsb_en_sync.oclk_i  = L_clk_i;
  assign \fsb_en_sync.z.bss.iclk_data_i  = R_en_i;
  assign \fsb_en_sync.z.bss.oclk_data_o  = \fsb_en_sync.z.bss.bsg_SYNC_2_r ;
  assign \fsb_en_sync.z.bss.oclk_i  = L_clk_i;
  assign \l2r_fifo.MSYNC_1r1w.r_addr_i  = \l2r_fifo.bapg_rd.w_ptr_r [0];
  assign \l2r_fifo.MSYNC_1r1w.r_data_o  = R_data_o;
  assign \l2r_fifo.MSYNC_1r1w.r_v_i  = R_v_o;
  assign \l2r_fifo.MSYNC_1r1w.synth.r_addr_i  = \l2r_fifo.bapg_rd.w_ptr_r [0];
  assign \l2r_fifo.MSYNC_1r1w.synth.r_data_o  = R_data_o;
  assign \l2r_fifo.MSYNC_1r1w.synth.r_v_i  = R_v_o;
  assign \l2r_fifo.MSYNC_1r1w.synth.unused0  = L_reset_i;
  assign \l2r_fifo.MSYNC_1r1w.synth.unused1  = R_v_o;
  assign \l2r_fifo.MSYNC_1r1w.synth.w_addr_i  = \l2r_fifo.bapg_wr.w_ptr_r [0];
  assign \l2r_fifo.MSYNC_1r1w.synth.w_clk_i  = L_clk_i;
  assign \l2r_fifo.MSYNC_1r1w.synth.w_data_i  = L_data_i;
  assign \l2r_fifo.MSYNC_1r1w.synth.w_reset_i  = L_reset_i;
  assign \l2r_fifo.MSYNC_1r1w.synth.w_v_i  = \l2r_fifo.bapg_wr.w_inc_i ;
  assign \l2r_fifo.MSYNC_1r1w.w_addr_i  = \l2r_fifo.bapg_wr.w_ptr_r [0];
  assign \l2r_fifo.MSYNC_1r1w.w_clk_i  = L_clk_i;
  assign \l2r_fifo.MSYNC_1r1w.w_data_i  = L_data_i;
  assign \l2r_fifo.MSYNC_1r1w.w_reset_i  = L_reset_i;
  assign \l2r_fifo.MSYNC_1r1w.w_v_i  = \l2r_fifo.bapg_wr.w_inc_i ;
  assign \l2r_fifo.bapg_rd.ptr_sync.iclk_data_o  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.bapg_rd.ptr_sync.iclk_i  = R_clk_i;
  assign \l2r_fifo.bapg_rd.ptr_sync.iclk_reset_i  = R_reset_i;
  assign \l2r_fifo.bapg_rd.ptr_sync.oclk_data_o  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.bapg_rd.ptr_sync.oclk_i  = L_clk_i;
  assign \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_data_o  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_i  = R_clk_i;
  assign \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_reset_i  = R_reset_i;
  assign \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.oclk_data_o  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.oclk_i  = L_clk_i;
  assign \l2r_fifo.bapg_rd.r_clk_i  = L_clk_i;
  assign \l2r_fifo.bapg_rd.w_clk_i  = R_clk_i;
  assign \l2r_fifo.bapg_rd.w_inc_i  = R_yumi_i;
  assign \l2r_fifo.bapg_rd.w_ptr_binary_r_o  = { 1'hx, \l2r_fifo.bapg_rd.w_ptr_r [0] };
  assign \l2r_fifo.bapg_rd.w_ptr_gray_r  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.bapg_rd.w_ptr_gray_r_o  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.bapg_rd.w_ptr_gray_r_rsync  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.bapg_rd.w_ptr_gray_r_rsync_o  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.bapg_rd.w_ptr_p1_r [1] = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  assign \l2r_fifo.bapg_rd.w_ptr_r [1] = 1'hx;
  assign \l2r_fifo.bapg_rd.w_reset_i  = R_reset_i;
  assign \l2r_fifo.bapg_wr.ptr_sync.iclk_data_o  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.bapg_wr.ptr_sync.iclk_i  = L_clk_i;
  assign \l2r_fifo.bapg_wr.ptr_sync.iclk_reset_i  = L_reset_i;
  assign \l2r_fifo.bapg_wr.ptr_sync.oclk_data_o  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.bapg_wr.ptr_sync.oclk_i  = R_clk_i;
  assign \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_data_o  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_i  = L_clk_i;
  assign \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_reset_i  = L_reset_i;
  assign \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.oclk_data_o  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.oclk_i  = R_clk_i;
  assign \l2r_fifo.bapg_wr.r_clk_i  = R_clk_i;
  assign \l2r_fifo.bapg_wr.w_clk_i  = L_clk_i;
  assign \l2r_fifo.bapg_wr.w_ptr_binary_r_o  = { 1'hx, \l2r_fifo.bapg_wr.w_ptr_r [0] };
  assign \l2r_fifo.bapg_wr.w_ptr_gray_r  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.bapg_wr.w_ptr_gray_r_o  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.bapg_wr.w_ptr_gray_r_rsync  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.bapg_wr.w_ptr_gray_r_rsync_o  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.bapg_wr.w_ptr_p1_r [1] = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  assign \l2r_fifo.bapg_wr.w_ptr_r [1] = 1'hx;
  assign \l2r_fifo.bapg_wr.w_reset_i  = L_reset_i;
  assign \l2r_fifo.r_clk_i  = R_clk_i;
  assign \l2r_fifo.r_data_o  = R_data_o;
  assign \l2r_fifo.r_data_o_tmp  = R_data_o;
  assign \l2r_fifo.r_deq_i  = R_yumi_i;
  assign \l2r_fifo.r_ptr_binary_r  = { 1'hx, \l2r_fifo.bapg_rd.w_ptr_r [0] };
  assign \l2r_fifo.r_ptr_gray_r  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.r_ptr_gray_r_wsync  = \l2r_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.r_reset_i  = R_reset_i;
  assign \l2r_fifo.r_valid_o  = R_v_o;
  assign \l2r_fifo.r_valid_o_tmp  = R_v_o;
  assign \l2r_fifo.w_clk_i  = L_clk_i;
  assign \l2r_fifo.w_data_i  = L_data_i;
  assign \l2r_fifo.w_enq_i  = \l2r_fifo.bapg_wr.w_inc_i ;
  assign \l2r_fifo.w_ptr_binary_r  = { 1'hx, \l2r_fifo.bapg_wr.w_ptr_r [0] };
  assign \l2r_fifo.w_ptr_gray_r  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \l2r_fifo.w_ptr_gray_r_rsync  = \l2r_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \l2r_fifo.w_reset_i  = L_reset_i;
  assign \r2l_fifo.MSYNC_1r1w.r_addr_i  = \r2l_fifo.bapg_rd.w_ptr_r [0];
  assign \r2l_fifo.MSYNC_1r1w.r_data_o  = L_data_o;
  assign \r2l_fifo.MSYNC_1r1w.r_v_i  = L_v_o;
  assign \r2l_fifo.MSYNC_1r1w.synth.r_addr_i  = \r2l_fifo.bapg_rd.w_ptr_r [0];
  assign \r2l_fifo.MSYNC_1r1w.synth.r_data_o  = L_data_o;
  assign \r2l_fifo.MSYNC_1r1w.synth.r_v_i  = L_v_o;
  assign \r2l_fifo.MSYNC_1r1w.synth.unused0  = R_reset_i;
  assign \r2l_fifo.MSYNC_1r1w.synth.unused1  = L_v_o;
  assign \r2l_fifo.MSYNC_1r1w.synth.w_addr_i  = \r2l_fifo.bapg_wr.w_ptr_r [0];
  assign \r2l_fifo.MSYNC_1r1w.synth.w_clk_i  = R_clk_i;
  assign \r2l_fifo.MSYNC_1r1w.synth.w_data_i  = R_data_i;
  assign \r2l_fifo.MSYNC_1r1w.synth.w_reset_i  = R_reset_i;
  assign \r2l_fifo.MSYNC_1r1w.synth.w_v_i  = \r2l_fifo.bapg_wr.w_inc_i ;
  assign \r2l_fifo.MSYNC_1r1w.w_addr_i  = \r2l_fifo.bapg_wr.w_ptr_r [0];
  assign \r2l_fifo.MSYNC_1r1w.w_clk_i  = R_clk_i;
  assign \r2l_fifo.MSYNC_1r1w.w_data_i  = R_data_i;
  assign \r2l_fifo.MSYNC_1r1w.w_reset_i  = R_reset_i;
  assign \r2l_fifo.MSYNC_1r1w.w_v_i  = \r2l_fifo.bapg_wr.w_inc_i ;
  assign \r2l_fifo.bapg_rd.ptr_sync.iclk_data_o  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.bapg_rd.ptr_sync.iclk_i  = L_clk_i;
  assign \r2l_fifo.bapg_rd.ptr_sync.iclk_reset_i  = L_reset_i;
  assign \r2l_fifo.bapg_rd.ptr_sync.oclk_data_o  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.bapg_rd.ptr_sync.oclk_i  = R_clk_i;
  assign \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_data_o  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_i  = L_clk_i;
  assign \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.iclk_reset_i  = L_reset_i;
  assign \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.oclk_data_o  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.oclk_i  = R_clk_i;
  assign \r2l_fifo.bapg_rd.r_clk_i  = R_clk_i;
  assign \r2l_fifo.bapg_rd.w_clk_i  = L_clk_i;
  assign \r2l_fifo.bapg_rd.w_ptr_binary_r_o  = { 1'hx, \r2l_fifo.bapg_rd.w_ptr_r [0] };
  assign \r2l_fifo.bapg_rd.w_ptr_gray_r  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.bapg_rd.w_ptr_gray_r_o  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.bapg_rd.w_ptr_gray_r_rsync  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.bapg_rd.w_ptr_gray_r_rsync_o  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.bapg_rd.w_ptr_p1_r [1] = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  assign \r2l_fifo.bapg_rd.w_ptr_r [1] = 1'hx;
  assign \r2l_fifo.bapg_rd.w_reset_i  = L_reset_i;
  assign \r2l_fifo.bapg_wr.ptr_sync.iclk_data_o  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.bapg_wr.ptr_sync.iclk_i  = R_clk_i;
  assign \r2l_fifo.bapg_wr.ptr_sync.iclk_reset_i  = R_reset_i;
  assign \r2l_fifo.bapg_wr.ptr_sync.oclk_data_o  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.bapg_wr.ptr_sync.oclk_i  = L_clk_i;
  assign \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_data_o  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_i  = R_clk_i;
  assign \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.iclk_reset_i  = R_reset_i;
  assign \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.oclk_data_o  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.oclk_i  = L_clk_i;
  assign \r2l_fifo.bapg_wr.r_clk_i  = L_clk_i;
  assign \r2l_fifo.bapg_wr.w_clk_i  = R_clk_i;
  assign \r2l_fifo.bapg_wr.w_ptr_binary_r_o  = { 1'hx, \r2l_fifo.bapg_wr.w_ptr_r [0] };
  assign \r2l_fifo.bapg_wr.w_ptr_gray_r  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.bapg_wr.w_ptr_gray_r_o  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.bapg_wr.w_ptr_gray_r_rsync  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.bapg_wr.w_ptr_gray_r_rsync_o  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.bapg_wr.w_ptr_p1_r [1] = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  assign \r2l_fifo.bapg_wr.w_ptr_r [1] = 1'hx;
  assign \r2l_fifo.bapg_wr.w_reset_i  = R_reset_i;
  assign \r2l_fifo.r_clk_i  = L_clk_i;
  assign \r2l_fifo.r_data_o  = L_data_o;
  assign \r2l_fifo.r_data_o_tmp  = L_data_o;
  assign \r2l_fifo.r_deq_i  = \r2l_fifo.bapg_rd.w_inc_i ;
  assign \r2l_fifo.r_ptr_binary_r  = { 1'hx, \r2l_fifo.bapg_rd.w_ptr_r [0] };
  assign \r2l_fifo.r_ptr_gray_r  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.r_ptr_gray_r_wsync  = \r2l_fifo.bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.r_reset_i  = L_reset_i;
  assign \r2l_fifo.r_valid_o  = L_v_o;
  assign \r2l_fifo.r_valid_o_tmp  = L_v_o;
  assign \r2l_fifo.w_clk_i  = R_clk_i;
  assign \r2l_fifo.w_data_i  = R_data_i;
  assign \r2l_fifo.w_enq_i  = \r2l_fifo.bapg_wr.w_inc_i ;
  assign \r2l_fifo.w_ptr_binary_r  = { 1'hx, \r2l_fifo.bapg_wr.w_ptr_r [0] };
  assign \r2l_fifo.w_ptr_gray_r  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \r2l_fifo.w_ptr_gray_r_rsync  = \r2l_fifo.bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \r2l_fifo.w_reset_i  = R_reset_i;
endmodule
