module bsg_arb_fixed(ready_i, reqs_i, grants_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire [15:0] \enc.i ;
  wire [15:0] \enc.nw1.scan.i ;
  wire [15:0] \enc.nw1.scan.o ;
  wire [15:0] \enc.nw1.scan.scanN.row[0].fill ;
  wire [15:0] \enc.nw1.scan.scanN.row[0].shifted ;
  wire [15:0] \enc.nw1.scan.scanN.row[1].fill ;
  wire [15:0] \enc.nw1.scan.scanN.row[1].shifted ;
  wire [15:0] \enc.nw1.scan.scanN.row[2].fill ;
  wire [15:0] \enc.nw1.scan.scanN.row[2].shifted ;
  wire [15:0] \enc.nw1.scan.scanN.row[3].fill ;
  wire [15:0] \enc.nw1.scan.scanN.row[3].shifted ;
  wire [79:0] \enc.nw1.scan.t ;
  wire [15:0] \enc.o ;
  wire [15:0] \enc.scan_lo ;
  wire \enc.v_o ;
  output [15:0] grants_o;
  wire [15:0] grants_o;
  wire [15:0] grants_unmasked_lo;
  input ready_i;
  wire ready_i;
  input [15:0] reqs_i;
  wire [15:0] reqs_i;
  assign _006_ = ~(reqs_i[1] | reqs_i[0]);
  assign _007_ = reqs_i[3] | reqs_i[2];
  assign _008_ = _006_ & ~(_007_);
  assign _009_ = reqs_i[5] | reqs_i[4];
  assign _010_ = reqs_i[7] | reqs_i[6];
  assign _011_ = _010_ | _009_;
  assign _012_ = _008_ & ~(_011_);
  assign _013_ = reqs_i[9] | reqs_i[8];
  assign _014_ = reqs_i[11] | reqs_i[10];
  assign _015_ = _014_ | _013_;
  assign _016_ = reqs_i[13] | reqs_i[12];
  assign _017_ = reqs_i[14] | reqs_i[15];
  assign _018_ = _017_ | _016_;
  assign _019_ = ~(_018_ | _015_);
  assign _020_ = ~(_019_ & _012_);
  assign _021_ = ~(reqs_i[2] | reqs_i[1]);
  assign _022_ = reqs_i[4] | reqs_i[3];
  assign _023_ = _021_ & ~(_022_);
  assign _024_ = reqs_i[6] | reqs_i[5];
  assign _025_ = reqs_i[8] | reqs_i[7];
  assign _026_ = _025_ | _024_;
  assign _027_ = _023_ & ~(_026_);
  assign _028_ = reqs_i[10] | reqs_i[9];
  assign _029_ = reqs_i[12] | reqs_i[11];
  assign _030_ = _029_ | _028_;
  assign _031_ = reqs_i[14] | reqs_i[13];
  assign _032_ = _031_ | reqs_i[15];
  assign _033_ = _032_ | _030_;
  assign _034_ = _027_ & ~(_033_);
  assign _035_ = ~(_034_ & _020_);
  assign grants_o[0] = ready_i & ~(_035_);
  assign _036_ = ~(_009_ | _007_);
  assign _037_ = _013_ | _010_;
  assign _038_ = _036_ & ~(_037_);
  assign _039_ = _016_ | _014_;
  assign _040_ = _039_ | _017_;
  assign _041_ = _038_ & ~(_040_);
  assign _042_ = _034_ | ~(_041_);
  assign grants_o[1] = ready_i & ~(_042_);
  assign _043_ = ~(_024_ | _022_);
  assign _044_ = _028_ | _025_;
  assign _045_ = _043_ & ~(_044_);
  assign _046_ = _031_ | _029_;
  assign _047_ = _046_ | reqs_i[15];
  assign _048_ = _045_ & ~(_047_);
  assign _049_ = _041_ | ~(_048_);
  assign grants_o[2] = ready_i & ~(_049_);
  assign _050_ = _015_ | _011_;
  assign _051_ = ~(_050_ | _018_);
  assign _052_ = _048_ | ~(_051_);
  assign grants_o[3] = ready_i & ~(_052_);
  assign _053_ = _030_ | _026_;
  assign _054_ = ~(_053_ | _032_);
  assign _055_ = _051_ | ~(_054_);
  assign grants_o[4] = ready_i & ~(_055_);
  assign _056_ = _039_ | _037_;
  assign _057_ = ~(_056_ | _017_);
  assign _058_ = _054_ | ~(_057_);
  assign grants_o[5] = ready_i & ~(_058_);
  assign _059_ = _046_ | _044_;
  assign _060_ = ~(_059_ | reqs_i[15]);
  assign _061_ = _057_ | ~(_060_);
  assign grants_o[6] = ready_i & ~(_061_);
  assign _062_ = _060_ | ~(_019_);
  assign grants_o[7] = ready_i & ~(_062_);
  assign _063_ = _033_ | _019_;
  assign grants_o[8] = ready_i & ~(_063_);
  assign _000_ = _040_ | ~(_033_);
  assign grants_o[9] = ready_i & ~(_000_);
  assign _001_ = _047_ | ~(_040_);
  assign grants_o[10] = ready_i & ~(_001_);
  assign _002_ = _018_ | ~(_047_);
  assign grants_o[11] = ready_i & ~(_002_);
  assign _003_ = _032_ | ~(_018_);
  assign grants_o[12] = ready_i & ~(_003_);
  assign _004_ = _017_ | ~(_032_);
  assign grants_o[13] = ready_i & ~(_004_);
  assign _005_ = reqs_i[15] | ~(reqs_i[14]);
  assign grants_o[14] = ready_i & ~(_005_);
  assign grants_o[15] = ready_i & reqs_i[15];
  assign \enc.i  = reqs_i;
  assign \enc.nw1.scan.i  = reqs_i;
  assign \enc.nw1.scan.o [15] = reqs_i[15];
  assign \enc.nw1.scan.scanN.row[0].fill  = 16'h0000;
  assign \enc.nw1.scan.scanN.row[0].shifted  = { 1'h0, reqs_i[15:1] };
  assign \enc.nw1.scan.scanN.row[1].fill  = 16'h0000;
  assign \enc.nw1.scan.scanN.row[1].shifted [15:12] = { 2'h0, reqs_i[15], \enc.nw1.scan.o [14] };
  assign \enc.nw1.scan.scanN.row[2].fill  = 16'h0000;
  assign \enc.nw1.scan.scanN.row[2].shifted [15:8] = { 4'h0, reqs_i[15], \enc.nw1.scan.o [14:12] };
  assign \enc.nw1.scan.scanN.row[3].fill  = 16'h0000;
  assign \enc.nw1.scan.scanN.row[3].shifted  = { 8'h00, reqs_i[15], \enc.nw1.scan.o [14:8] };
  assign { \enc.nw1.scan.t [79:56], \enc.nw1.scan.t [47:36], \enc.nw1.scan.t [31:18], \enc.nw1.scan.t [15:0] } = { reqs_i[15], \enc.nw1.scan.o [14:0], reqs_i[15], \enc.nw1.scan.o [14:8], reqs_i[15], \enc.nw1.scan.o [14:12], \enc.nw1.scan.scanN.row[2].shifted [7:0], reqs_i[15], \enc.nw1.scan.o [14], \enc.nw1.scan.scanN.row[1].shifted [11:0], reqs_i };
  assign \enc.o [15] = reqs_i[15];
  assign \enc.scan_lo  = { reqs_i[15], \enc.nw1.scan.o [14:0] };
  assign \enc.v_o  = \enc.nw1.scan.o [0];
  assign grants_unmasked_lo = { reqs_i[15], \enc.o [14:0] };
endmodule
