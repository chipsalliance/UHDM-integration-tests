module bsg_less_than(a_i, b_i, o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  input [15:0] a_i;
  wire [15:0] a_i;
  input [15:0] b_i;
  wire [15:0] b_i;
  output o;
  wire o;
  assign _011_ = b_i[15] & ~(a_i[15]);
  assign _012_ = ~(b_i[15] ^ a_i[15]);
  assign _013_ = a_i[14] | ~(b_i[14]);
  assign _014_ = _012_ & ~(_013_);
  assign _015_ = _014_ | _011_;
  assign _016_ = b_i[14] ^ a_i[14];
  assign _017_ = _012_ & ~(_016_);
  assign _018_ = a_i[13] | ~(b_i[13]);
  assign _019_ = b_i[13] ^ a_i[13];
  assign _020_ = b_i[12] & ~(a_i[12]);
  assign _021_ = _020_ & ~(_019_);
  assign _022_ = _018_ & ~(_021_);
  assign _023_ = _017_ & ~(_022_);
  assign _024_ = _023_ | _015_;
  assign _025_ = b_i[12] ^ a_i[12];
  assign _026_ = _025_ | _019_;
  assign _027_ = _017_ & ~(_026_);
  assign _028_ = a_i[11] | ~(b_i[11]);
  assign _029_ = ~(b_i[11] ^ a_i[11]);
  assign _030_ = a_i[10] | ~(b_i[10]);
  assign _031_ = _029_ & ~(_030_);
  assign _032_ = _028_ & ~(_031_);
  assign _033_ = b_i[10] ^ a_i[10];
  assign _034_ = _033_ | ~(_029_);
  assign _035_ = a_i[9] | ~(b_i[9]);
  assign _036_ = b_i[9] ^ a_i[9];
  assign _037_ = b_i[8] & ~(a_i[8]);
  assign _038_ = _037_ & ~(_036_);
  assign _039_ = _038_ | ~(_035_);
  assign _040_ = _039_ & ~(_034_);
  assign _041_ = _032_ & ~(_040_);
  assign _042_ = _027_ & ~(_041_);
  assign _043_ = _042_ | _024_;
  assign _044_ = b_i[8] ^ a_i[8];
  assign _045_ = _044_ | _036_;
  assign _046_ = _045_ | _034_;
  assign _047_ = _027_ & ~(_046_);
  assign _048_ = a_i[7] | ~(b_i[7]);
  assign _049_ = ~(b_i[7] ^ a_i[7]);
  assign _050_ = a_i[6] | ~(b_i[6]);
  assign _051_ = _049_ & ~(_050_);
  assign _052_ = _048_ & ~(_051_);
  assign _053_ = b_i[6] ^ a_i[6];
  assign _054_ = _049_ & ~(_053_);
  assign _055_ = a_i[5] | ~(b_i[5]);
  assign _056_ = b_i[5] ^ a_i[5];
  assign _057_ = b_i[4] & ~(a_i[4]);
  assign _058_ = _057_ & ~(_056_);
  assign _059_ = _055_ & ~(_058_);
  assign _060_ = _054_ & ~(_059_);
  assign _061_ = _052_ & ~(_060_);
  assign _062_ = b_i[4] ^ a_i[4];
  assign _063_ = _062_ | _056_;
  assign _064_ = _063_ | ~(_054_);
  assign _065_ = a_i[3] | ~(b_i[3]);
  assign _066_ = ~(b_i[3] ^ a_i[3]);
  assign _067_ = a_i[2] | ~(b_i[2]);
  assign _068_ = _066_ & ~(_067_);
  assign _069_ = _065_ & ~(_068_);
  assign _070_ = b_i[2] ^ a_i[2];
  assign _071_ = _070_ | ~(_066_);
  assign _072_ = a_i[1] | ~(b_i[1]);
  assign _073_ = b_i[1] ^ a_i[1];
  assign _074_ = b_i[0] | ~(a_i[0]);
  assign _075_ = _074_ & ~(_073_);
  assign _076_ = _075_ | ~(_072_);
  assign _000_ = _076_ & ~(_071_);
  assign _001_ = _000_ | ~(_069_);
  assign _002_ = _001_ & ~(_064_);
  assign _003_ = _061_ & ~(_002_);
  assign _004_ = _047_ & ~(_003_);
  assign _005_ = _004_ | _043_;
  assign _006_ = b_i[0] ^ a_i[0];
  assign _007_ = _006_ | _073_;
  assign _008_ = _007_ | _071_;
  assign _009_ = _008_ | _064_;
  assign _010_ = _047_ & ~(_009_);
  assign o = _005_ & ~(_010_);
endmodule
