module bsg_mux_bitwise(data0_i, data1_i, sel_i, data_o);
  input [15:0] data0_i;
  wire [15:0] data0_i;
  input [15:0] data1_i;
  wire [15:0] data1_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire [15:0] \mux_segmented.data0_i ;
  wire [15:0] \mux_segmented.data1_i ;
  wire [15:0] \mux_segmented.data_o ;
  wire [15:0] \mux_segmented.sel_i ;
  input [15:0] sel_i;
  wire [15:0] sel_i;
  assign data_o[9] = sel_i[9] ? data1_i[9] : data0_i[9];
  assign data_o[8] = sel_i[8] ? data1_i[8] : data0_i[8];
  assign data_o[7] = sel_i[7] ? data1_i[7] : data0_i[7];
  assign data_o[6] = sel_i[6] ? data1_i[6] : data0_i[6];
  assign data_o[5] = sel_i[5] ? data1_i[5] : data0_i[5];
  assign data_o[4] = sel_i[4] ? data1_i[4] : data0_i[4];
  assign data_o[3] = sel_i[3] ? data1_i[3] : data0_i[3];
  assign data_o[2] = sel_i[2] ? data1_i[2] : data0_i[2];
  assign data_o[1] = sel_i[1] ? data1_i[1] : data0_i[1];
  assign data_o[0] = sel_i[0] ? data1_i[0] : data0_i[0];
  assign data_o[15] = sel_i[15] ? data1_i[15] : data0_i[15];
  assign data_o[14] = sel_i[14] ? data1_i[14] : data0_i[14];
  assign data_o[13] = sel_i[13] ? data1_i[13] : data0_i[13];
  assign data_o[12] = sel_i[12] ? data1_i[12] : data0_i[12];
  assign data_o[11] = sel_i[11] ? data1_i[11] : data0_i[11];
  assign data_o[10] = sel_i[10] ? data1_i[10] : data0_i[10];
  assign \mux_segmented.data0_i  = data0_i;
  assign \mux_segmented.data1_i  = data1_i;
  assign \mux_segmented.data_o  = data_o;
  assign \mux_segmented.sel_i  = sel_i;
endmodule
