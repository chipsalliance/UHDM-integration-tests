module bsg_flow_convert(v_i, fc_o, v_o, fc_i);
  input fc_i;
  wire fc_i;
  output fc_o;
  wire fc_o;
  input v_i;
  wire v_i;
  output v_o;
  wire v_o;
  assign fc_o = fc_i;
  assign v_o = v_i;
endmodule
