module bsg_channel_narrow(clk_i, reset_i, data_i, deque_o, data_o, deque_i);
  input clk_i;
  wire clk_i;
  wire count_n;
  reg count_r;
  wire [7:0] \data[0] ;
  wire [7:0] \data[1] ;
  input [15:0] data_i;
  wire [15:0] data_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  input deque_i;
  wire deque_i;
  output deque_o;
  wire deque_o;
  input reset_i;
  wire reset_i;
  assign data_o[0] = count_r ? data_i[8] : data_i[0];
  assign data_o[1] = count_r ? data_i[9] : data_i[1];
  assign data_o[2] = count_r ? data_i[10] : data_i[2];
  assign data_o[3] = count_r ? data_i[11] : data_i[3];
  assign data_o[4] = count_r ? data_i[12] : data_i[4];
  assign data_o[5] = count_r ? data_i[13] : data_i[5];
  assign data_o[6] = count_r ? data_i[14] : data_i[6];
  assign data_o[7] = count_r ? data_i[15] : data_i[7];
  assign count_n = deque_i ^ count_r;
  assign deque_o = deque_i & count_r;
  always @(posedge clk_i)
    if (reset_i) count_r <= 1'h0;
    else count_r <= count_n;
  assign \data[0]  = data_i[7:0];
  assign \data[1]  = data_i[15:8];
endmodule
