module dut (output int o);
  assign o = 1;
endmodule
