module top;
   int a = '0;
   int b = '1;
   int c = 'x;
   int d = 'z;
endmodule // top
