module bsg_buf_ctrl(i, o);
  input i;
  wire i;
  output [15:0] o;
  wire [15:0] o;
  assign o = { i, i, i, i, i, i, i, i, i, i, i, i, i, i, i, i };
endmodule
