module bsg_fpu_preprocess(a_i, zero_o, nan_o, sig_nan_o, infty_o, exp_zero_o, man_zero_o, denormal_o, sign_o, exp_o, man_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  input [15:0] a_i;
  wire [15:0] a_i;
  output denormal_o;
  wire denormal_o;
  output [4:0] exp_o;
  wire [4:0] exp_o;
  wire exp_zero;
  output exp_zero_o;
  wire exp_zero_o;
  output infty_o;
  wire infty_o;
  output [9:0] man_o;
  wire [9:0] man_o;
  output man_zero_o;
  wire man_zero_o;
  wire mantissa_zero;
  output nan_o;
  wire nan_o;
  output sig_nan_o;
  wire sig_nan_o;
  output sign_o;
  wire sign_o;
  output zero_o;
  wire zero_o;
  assign _00_ = ~(a_i[1] | a_i[0]);
  assign _01_ = a_i[3] | a_i[2];
  assign _02_ = _00_ & ~(_01_);
  assign _03_ = a_i[5] | a_i[4];
  assign _04_ = a_i[7] | a_i[6];
  assign _05_ = _04_ | _03_;
  assign _06_ = _02_ & ~(_05_);
  assign _07_ = a_i[9] | a_i[8];
  assign man_zero_o = _06_ & ~(_07_);
  assign _08_ = ~a_i[14];
  assign _09_ = a_i[11] | a_i[10];
  assign _10_ = a_i[13] | a_i[12];
  assign _11_ = _10_ | _09_;
  assign exp_zero_o = _08_ & ~(_11_);
  assign _12_ = ~exp_zero_o;
  assign zero_o = man_zero_o & ~(_12_);
  assign _13_ = ~(a_i[11] & a_i[10]);
  assign _14_ = ~(a_i[13] & a_i[12]);
  assign _15_ = _14_ | _13_;
  assign _16_ = _15_ | _08_;
  assign nan_o = ~(_16_ | man_zero_o);
  assign sig_nan_o = nan_o & ~(a_i[9]);
  assign infty_o = man_zero_o & ~(_16_);
  assign denormal_o = ~(_12_ | man_zero_o);
  assign exp_o = a_i[14:10];
  assign exp_zero = exp_zero_o;
  assign man_o = a_i[9:0];
  assign mantissa_zero = man_zero_o;
  assign sign_o = a_i[15];
endmodule
