module top(output int o);
   assign o = int'(50us);
endmodule
