module bsg_decode_with_v(i, v_i, o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire [3:0] \bd.i ;
  input [3:0] i;
  wire [3:0] i;
  output [15:0] o;
  wire [15:0] o;
  input v_i;
  wire v_i;
  assign _00_ = i[0] | i[1];
  assign _01_ = _00_ | i[2];
  assign _02_ = _01_ | i[3];
  assign o[0] = v_i & ~(_02_);
  assign _03_ = i[1] | ~(i[0]);
  assign _04_ = _03_ | i[2];
  assign _05_ = _04_ | i[3];
  assign o[1] = v_i & ~(_05_);
  assign _06_ = i[0] | ~(i[1]);
  assign _07_ = _06_ | i[2];
  assign _08_ = _07_ | i[3];
  assign o[2] = v_i & ~(_08_);
  assign _09_ = ~(i[0] & i[1]);
  assign _10_ = _09_ | i[2];
  assign _11_ = _10_ | i[3];
  assign o[3] = v_i & ~(_11_);
  assign _12_ = ~i[2];
  assign _13_ = _00_ | _12_;
  assign _14_ = _13_ | i[3];
  assign o[4] = v_i & ~(_14_);
  assign _15_ = _03_ | _12_;
  assign _16_ = _15_ | i[3];
  assign o[5] = v_i & ~(_16_);
  assign _17_ = _06_ | _12_;
  assign _18_ = _17_ | i[3];
  assign o[6] = v_i & ~(_18_);
  assign _19_ = _09_ | _12_;
  assign _20_ = _19_ | i[3];
  assign o[7] = v_i & ~(_20_);
  assign _21_ = ~i[3];
  assign _22_ = _01_ | _21_;
  assign o[8] = v_i & ~(_22_);
  assign _23_ = _04_ | _21_;
  assign o[9] = v_i & ~(_23_);
  assign _24_ = _07_ | _21_;
  assign o[10] = v_i & ~(_24_);
  assign _25_ = _10_ | _21_;
  assign o[11] = v_i & ~(_25_);
  assign _26_ = _13_ | _21_;
  assign o[12] = v_i & ~(_26_);
  assign _27_ = _15_ | _21_;
  assign o[13] = v_i & ~(_27_);
  assign _28_ = _17_ | _21_;
  assign o[14] = v_i & ~(_28_);
  assign _29_ = _19_ | _21_;
  assign o[15] = v_i & ~(_29_);
  assign \bd.i  = i;
endmodule
