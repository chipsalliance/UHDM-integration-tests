module bsg_imul_iterative(clk_i, reset_i, v_i, ready_o, opA_i, signed_opA_i, opB_i, signed_opB_i, gets_high_part_i, v_o, result_o, yumi_i);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire [5:0] _0746_;
  wire [5:0] _0747_;
  reg all_sh_lsb_zero_r;
  input clk_i;
  wire clk_i;
  reg [5:0] curr_state_r;
  input gets_high_part_i;
  wire gets_high_part_i;
  reg gets_high_part_r;
  wire latch_input;
  reg need_neg_result_r;
  input [31:0] opA_i;
  wire [31:0] opA_i;
  reg [31:0] opA_r;
  input [31:0] opB_i;
  wire [31:0] opB_i;
  reg [31:0] opB_r;
  output ready_o;
  wire ready_o;
  input reset_i;
  wire reset_i;
  output [31:0] result_o;
  wire [31:0] result_o;
  reg [31:0] result_r;
  reg [5:0] shift_counter_r;
  wire signed_opA;
  input signed_opA_i;
  wire signed_opA_i;
  reg signed_opA_r;
  wire signed_opB;
  input signed_opB_i;
  wire signed_opB_i;
  reg signed_opB_r;
  input v_i;
  wire v_i;
  output v_o;
  wire v_o;
  input yumi_i;
  wire yumi_i;
  assign _0746_[0] = ~shift_counter_r[0];
  assign _0039_ = need_neg_result_r & curr_state_r[1];
  assign _0040_ = opB_r[0] & curr_state_r[5];
  assign _0041_ = _0040_ | _0039_;
  assign _0042_ = curr_state_r[5] & ~(opB_r[0]);
  assign _0043_ = _0042_ | _0041_;
  assign _0044_ = ~gets_high_part_r;
  assign _0045_ = _0044_ & ~(_0039_);
  assign _0046_ = opB_r[0] | ~(curr_state_r[5]);
  assign _0047_ = _0045_ & ~(_0046_);
  assign _0007_ = _0043_ & ~(_0047_);
  assign _0048_ = curr_state_r[1] & ~(reset_i);
  assign _0049_ = reset_i | yumi_i;
  assign _0050_ = curr_state_r[4] & ~(_0049_);
  assign _0010_ = _0050_ | _0048_;
  assign latch_input = curr_state_r[0] & v_i;
  assign _0051_ = reset_i | v_i;
  assign _0052_ = curr_state_r[0] & ~(_0051_);
  assign _0053_ = _0052_ | reset_i;
  assign _0054_ = reset_i | ~(yumi_i);
  assign _0055_ = curr_state_r[4] & ~(_0054_);
  assign _0003_ = _0055_ | _0053_;
  assign _0056_ = curr_state_r[0] | curr_state_r[1];
  assign _0057_ = curr_state_r[2] | curr_state_r[3];
  assign _0058_ = _0057_ | _0056_;
  assign _0059_ = _0058_ | curr_state_r[4];
  assign _0060_ = curr_state_r[4] & ~(yumi_i);
  assign _0061_ = ~(_0060_ | curr_state_r[1]);
  assign _0062_ = ~(gets_high_part_r ^ shift_counter_r[0]);
  assign _0063_ = shift_counter_r[1] ^ gets_high_part_r;
  assign _0064_ = _0062_ & ~(_0063_);
  assign _0065_ = shift_counter_r[2] ^ gets_high_part_r;
  assign _0066_ = shift_counter_r[3] ^ gets_high_part_r;
  assign _0067_ = _0066_ | _0065_;
  assign _0068_ = _0064_ & ~(_0067_);
  assign _0069_ = shift_counter_r[4] ^ gets_high_part_r;
  assign _0070_ = ~(shift_counter_r[5] ^ gets_high_part_r);
  assign _0071_ = _0070_ | _0069_;
  assign _0072_ = _0068_ & ~(_0071_);
  assign _0073_ = curr_state_r[5] & ~(_0072_);
  assign _0074_ = _0073_ | curr_state_r[2];
  assign _0075_ = _0061_ & ~(_0074_);
  assign _0076_ = _0075_ & ~(latch_input);
  assign _0077_ = ~(curr_state_r[4] | curr_state_r[1]);
  assign _0078_ = curr_state_r[5] | curr_state_r[2];
  assign _0079_ = _0077_ & ~(_0078_);
  assign _0080_ = curr_state_r[0] | curr_state_r[3];
  assign _0081_ = _0079_ & ~(_0080_);
  assign _0082_ = _0081_ | _0076_;
  assign _0083_ = ~(_0074_ | curr_state_r[3]);
  assign _0084_ = _0083_ | _0081_;
  assign _0085_ = _0084_ | _0082_;
  assign _0086_ = ~curr_state_r[5];
  assign _0087_ = _0072_ & ~(_0086_);
  assign _0088_ = _0087_ | ~(_0061_);
  assign _0089_ = _0088_ & ~(_0081_);
  assign _0090_ = _0089_ | _0085_;
  assign _0091_ = _0059_ & ~(_0090_);
  assign _0008_ = _0091_ | reset_i;
  assign _0009_ = latch_input | reset_i;
  assign _0006_ = latch_input | curr_state_r[5];
  assign _0092_ = signed_opB_r & curr_state_r[2];
  assign _0093_ = _0092_ | latch_input;
  assign _0005_ = _0093_ | curr_state_r[5];
  assign _0094_ = curr_state_r[2] & ~(reset_i);
  assign _0095_ = _0072_ | reset_i;
  assign _0096_ = curr_state_r[5] & ~(_0095_);
  assign _0011_ = _0096_ | _0094_;
  assign _0097_ = curr_state_r[5] & ~(gets_high_part_r);
  assign _0098_ = _0097_ | latch_input;
  assign _0099_ = signed_opA_r & curr_state_r[3];
  assign _0004_ = _0099_ | _0098_;
  assign _0100_ = ~_0040_;
  assign _0101_ = ~(result_r[0] ^ curr_state_r[1]);
  assign _0102_ = curr_state_r[2] ? opB_r[0] : _0101_;
  assign _0103_ = curr_state_r[3] ? opA_r[0] : _0102_;
  assign _0104_ = _0057_ | curr_state_r[1];
  assign _0105_ = ~(_0104_ | opA_r[0]);
  assign _0106_ = ~(_0105_ ^ _0103_);
  assign _0107_ = ~_0106_;
  assign _0108_ = ~opA_r[1];
  assign _0109_ = ~opB_r[1];
  assign _0110_ = result_r[1] ^ curr_state_r[1];
  assign _0111_ = curr_state_r[2] ? _0109_ : _0110_;
  assign _0112_ = curr_state_r[3] ? _0108_ : _0111_;
  assign _0113_ = _0104_ | _0108_;
  assign _0114_ = ~(_0113_ ^ _0112_);
  assign _0115_ = _0105_ | _0103_;
  assign _0116_ = ~(_0115_ ^ _0114_);
  assign _0117_ = gets_high_part_r ? _0116_ : _0107_;
  assign _0118_ = _0040_ ? _0117_ : result_r[1];
  assign _0119_ = ~result_r[0];
  assign _0120_ = gets_high_part_r & ~(all_sh_lsb_zero_r);
  assign _0121_ = _0120_ ? _0119_ : _0107_;
  assign _0712_ = _0039_ ? _0121_ : _0118_;
  assign _0122_ = ~(result_r[2] ^ curr_state_r[1]);
  assign _0123_ = curr_state_r[2] ? opB_r[2] : _0122_;
  assign _0124_ = curr_state_r[3] ? opA_r[2] : _0123_;
  assign _0125_ = _0104_ | ~(opA_r[2]);
  assign _0126_ = ~(_0125_ ^ _0124_);
  assign _0127_ = _0112_ & ~(_0113_);
  assign _0128_ = _0114_ & ~(_0115_);
  assign _0129_ = _0128_ | _0127_;
  assign _0130_ = ~(_0129_ ^ _0126_);
  assign _0131_ = gets_high_part_r ? _0130_ : _0116_;
  assign _0132_ = _0040_ ? _0131_ : result_r[2];
  assign _0133_ = ~result_r[1];
  assign _0134_ = _0120_ ? _0133_ : _0116_;
  assign _0723_ = _0039_ ? _0134_ : _0132_;
  assign _0135_ = ~(result_r[3] ^ curr_state_r[1]);
  assign _0136_ = curr_state_r[2] ? opB_r[3] : _0135_;
  assign _0137_ = curr_state_r[3] ? opA_r[3] : _0136_;
  assign _0138_ = _0104_ | ~(opA_r[3]);
  assign _0139_ = ~(_0138_ ^ _0137_);
  assign _0140_ = _0125_ | _0124_;
  assign _0141_ = _0129_ & ~(_0126_);
  assign _0142_ = _0140_ & ~(_0141_);
  assign _0143_ = _0142_ ^ _0139_;
  assign _0144_ = gets_high_part_r ? _0143_ : _0130_;
  assign _0145_ = _0040_ ? _0144_ : result_r[3];
  assign _0146_ = ~result_r[2];
  assign _0147_ = _0120_ ? _0146_ : _0130_;
  assign _0734_ = _0039_ ? _0147_ : _0145_;
  assign _0148_ = ~(result_r[4] ^ curr_state_r[1]);
  assign _0149_ = curr_state_r[2] ? opB_r[4] : _0148_;
  assign _0150_ = curr_state_r[3] ? opA_r[4] : _0149_;
  assign _0151_ = _0104_ | ~(opA_r[4]);
  assign _0152_ = ~(_0151_ ^ _0150_);
  assign _0153_ = ~(_0138_ | _0137_);
  assign _0154_ = ~(_0140_ | _0139_);
  assign _0155_ = _0154_ | _0153_;
  assign _0156_ = _0139_ | _0126_;
  assign _0157_ = _0129_ & ~(_0156_);
  assign _0158_ = _0157_ | _0155_;
  assign _0159_ = ~(_0158_ ^ _0152_);
  assign _0160_ = gets_high_part_r ? _0159_ : _0143_;
  assign _0161_ = _0040_ ? _0160_ : result_r[4];
  assign _0162_ = ~result_r[3];
  assign _0163_ = _0120_ ? _0162_ : _0143_;
  assign _0737_ = _0039_ ? _0163_ : _0161_;
  assign _0164_ = ~(result_r[5] ^ curr_state_r[1]);
  assign _0165_ = curr_state_r[2] ? opB_r[5] : _0164_;
  assign _0166_ = curr_state_r[3] ? opA_r[5] : _0165_;
  assign _0167_ = _0104_ | ~(opA_r[5]);
  assign _0168_ = ~(_0167_ ^ _0166_);
  assign _0169_ = _0151_ | _0150_;
  assign _0170_ = _0158_ & ~(_0152_);
  assign _0171_ = _0169_ & ~(_0170_);
  assign _0172_ = _0171_ ^ _0168_;
  assign _0173_ = gets_high_part_r ? _0172_ : _0159_;
  assign _0174_ = _0040_ ? _0173_ : result_r[5];
  assign _0175_ = ~result_r[4];
  assign _0176_ = _0120_ ? _0175_ : _0159_;
  assign _0738_ = _0039_ ? _0176_ : _0174_;
  assign _0177_ = ~(result_r[6] ^ curr_state_r[1]);
  assign _0178_ = curr_state_r[2] ? opB_r[6] : _0177_;
  assign _0179_ = curr_state_r[3] ? opA_r[6] : _0178_;
  assign _0180_ = _0104_ | ~(opA_r[6]);
  assign _0181_ = ~(_0180_ ^ _0179_);
  assign _0182_ = ~(_0167_ | _0166_);
  assign _0183_ = ~(_0169_ | _0168_);
  assign _0184_ = _0183_ | _0182_;
  assign _0185_ = _0168_ | _0152_;
  assign _0186_ = _0185_ | ~(_0158_);
  assign _0187_ = _0186_ & ~(_0184_);
  assign _0188_ = _0187_ ^ _0181_;
  assign _0189_ = gets_high_part_r ? _0188_ : _0172_;
  assign _0190_ = _0040_ ? _0189_ : result_r[6];
  assign _0191_ = ~result_r[5];
  assign _0192_ = _0120_ ? _0191_ : _0172_;
  assign _0739_ = _0039_ ? _0192_ : _0190_;
  assign _0193_ = ~(result_r[7] ^ curr_state_r[1]);
  assign _0194_ = curr_state_r[2] ? opB_r[7] : _0193_;
  assign _0195_ = curr_state_r[3] ? opA_r[7] : _0194_;
  assign _0196_ = _0104_ | ~(opA_r[7]);
  assign _0197_ = ~(_0196_ ^ _0195_);
  assign _0198_ = _0180_ | _0179_;
  assign _0199_ = ~(_0187_ | _0181_);
  assign _0200_ = _0198_ & ~(_0199_);
  assign _0201_ = _0200_ ^ _0197_;
  assign _0202_ = gets_high_part_r ? _0201_ : _0188_;
  assign _0203_ = _0040_ ? _0202_ : result_r[7];
  assign _0204_ = ~result_r[6];
  assign _0205_ = _0120_ ? _0204_ : _0188_;
  assign _0740_ = _0039_ ? _0205_ : _0203_;
  assign _0206_ = ~(result_r[8] ^ curr_state_r[1]);
  assign _0207_ = curr_state_r[2] ? opB_r[8] : _0206_;
  assign _0208_ = curr_state_r[3] ? opA_r[8] : _0207_;
  assign _0209_ = _0104_ | ~(opA_r[8]);
  assign _0210_ = ~(_0209_ ^ _0208_);
  assign _0211_ = ~(_0196_ | _0195_);
  assign _0212_ = ~(_0198_ | _0197_);
  assign _0213_ = _0212_ | _0211_;
  assign _0214_ = _0197_ | _0181_;
  assign _0215_ = _0184_ & ~(_0214_);
  assign _0216_ = _0215_ | _0213_;
  assign _0217_ = _0214_ | _0185_;
  assign _0218_ = _0158_ & ~(_0217_);
  assign _0219_ = _0218_ | _0216_;
  assign _0220_ = ~(_0219_ ^ _0210_);
  assign _0221_ = gets_high_part_r ? _0220_ : _0201_;
  assign _0222_ = _0040_ ? _0221_ : result_r[8];
  assign _0223_ = ~result_r[7];
  assign _0224_ = _0120_ ? _0223_ : _0201_;
  assign _0741_ = _0039_ ? _0224_ : _0222_;
  assign _0225_ = ~(result_r[9] ^ curr_state_r[1]);
  assign _0226_ = curr_state_r[2] ? opB_r[9] : _0225_;
  assign _0227_ = curr_state_r[3] ? opA_r[9] : _0226_;
  assign _0228_ = _0104_ | ~(opA_r[9]);
  assign _0229_ = ~(_0228_ ^ _0227_);
  assign _0230_ = _0209_ | _0208_;
  assign _0231_ = _0219_ & ~(_0210_);
  assign _0232_ = _0230_ & ~(_0231_);
  assign _0233_ = _0232_ ^ _0229_;
  assign _0234_ = gets_high_part_r ? _0233_ : _0220_;
  assign _0235_ = _0040_ ? _0234_ : result_r[9];
  assign _0236_ = ~result_r[8];
  assign _0237_ = _0120_ ? _0236_ : _0220_;
  assign _0742_ = _0039_ ? _0237_ : _0235_;
  assign _0238_ = ~(result_r[10] ^ curr_state_r[1]);
  assign _0239_ = curr_state_r[2] ? opB_r[10] : _0238_;
  assign _0240_ = curr_state_r[3] ? opA_r[10] : _0239_;
  assign _0241_ = _0104_ | ~(opA_r[10]);
  assign _0242_ = ~(_0241_ ^ _0240_);
  assign _0243_ = ~(_0228_ | _0227_);
  assign _0244_ = ~(_0230_ | _0229_);
  assign _0245_ = _0244_ | _0243_;
  assign _0246_ = _0229_ | _0210_;
  assign _0247_ = _0246_ | ~(_0219_);
  assign _0248_ = _0247_ & ~(_0245_);
  assign _0249_ = _0248_ ^ _0242_;
  assign _0250_ = gets_high_part_r ? _0249_ : _0233_;
  assign _0251_ = _0040_ ? _0250_ : result_r[10];
  assign _0252_ = ~result_r[9];
  assign _0253_ = _0120_ ? _0252_ : _0233_;
  assign _0743_ = _0039_ ? _0253_ : _0251_;
  assign _0254_ = ~(result_r[11] ^ curr_state_r[1]);
  assign _0255_ = curr_state_r[2] ? opB_r[11] : _0254_;
  assign _0256_ = curr_state_r[3] ? opA_r[11] : _0255_;
  assign _0257_ = _0104_ | ~(opA_r[11]);
  assign _0258_ = ~(_0257_ ^ _0256_);
  assign _0259_ = _0241_ | _0240_;
  assign _0260_ = ~(_0248_ | _0242_);
  assign _0261_ = _0259_ & ~(_0260_);
  assign _0262_ = _0261_ ^ _0258_;
  assign _0263_ = gets_high_part_r ? _0262_ : _0249_;
  assign _0264_ = _0040_ ? _0263_ : result_r[11];
  assign _0265_ = ~result_r[10];
  assign _0266_ = _0120_ ? _0265_ : _0249_;
  assign _0713_ = _0039_ ? _0266_ : _0264_;
  assign _0267_ = ~(result_r[12] ^ curr_state_r[1]);
  assign _0268_ = curr_state_r[2] ? opB_r[12] : _0267_;
  assign _0269_ = curr_state_r[3] ? opA_r[12] : _0268_;
  assign _0270_ = _0104_ | ~(opA_r[12]);
  assign _0271_ = ~(_0270_ ^ _0269_);
  assign _0272_ = ~(_0257_ | _0256_);
  assign _0273_ = ~(_0259_ | _0258_);
  assign _0274_ = _0273_ | _0272_;
  assign _0275_ = _0258_ | _0242_;
  assign _0276_ = _0245_ & ~(_0275_);
  assign _0277_ = _0276_ | _0274_;
  assign _0278_ = _0275_ | _0246_;
  assign _0279_ = _0219_ & ~(_0278_);
  assign _0280_ = ~(_0279_ | _0277_);
  assign _0281_ = _0280_ ^ _0271_;
  assign _0282_ = gets_high_part_r ? _0281_ : _0262_;
  assign _0283_ = _0040_ ? _0282_ : result_r[12];
  assign _0284_ = ~result_r[11];
  assign _0285_ = _0120_ ? _0284_ : _0262_;
  assign _0714_ = _0039_ ? _0285_ : _0283_;
  assign _0286_ = ~(result_r[13] ^ curr_state_r[1]);
  assign _0287_ = curr_state_r[2] ? opB_r[13] : _0286_;
  assign _0288_ = curr_state_r[3] ? opA_r[13] : _0287_;
  assign _0289_ = _0104_ | ~(opA_r[13]);
  assign _0290_ = ~(_0289_ ^ _0288_);
  assign _0291_ = _0270_ | _0269_;
  assign _0292_ = ~(_0280_ | _0271_);
  assign _0293_ = _0291_ & ~(_0292_);
  assign _0294_ = _0293_ ^ _0290_;
  assign _0295_ = gets_high_part_r ? _0294_ : _0281_;
  assign _0296_ = _0040_ ? _0295_ : result_r[13];
  assign _0297_ = ~result_r[12];
  assign _0298_ = _0120_ ? _0297_ : _0281_;
  assign _0715_ = _0039_ ? _0298_ : _0296_;
  assign _0299_ = ~(result_r[14] ^ curr_state_r[1]);
  assign _0300_ = curr_state_r[2] ? opB_r[14] : _0299_;
  assign _0301_ = curr_state_r[3] ? opA_r[14] : _0300_;
  assign _0302_ = _0104_ | ~(opA_r[14]);
  assign _0303_ = ~(_0302_ ^ _0301_);
  assign _0304_ = ~(_0289_ | _0288_);
  assign _0305_ = ~(_0291_ | _0290_);
  assign _0306_ = _0305_ | _0304_;
  assign _0307_ = _0290_ | _0271_;
  assign _0308_ = _0307_ | _0280_;
  assign _0309_ = _0308_ & ~(_0306_);
  assign _0310_ = _0309_ ^ _0303_;
  assign _0311_ = gets_high_part_r ? _0310_ : _0294_;
  assign _0312_ = _0040_ ? _0311_ : result_r[14];
  assign _0313_ = ~result_r[13];
  assign _0314_ = _0120_ ? _0313_ : _0294_;
  assign _0716_ = _0039_ ? _0314_ : _0312_;
  assign _0315_ = ~(result_r[15] ^ curr_state_r[1]);
  assign _0316_ = curr_state_r[2] ? opB_r[15] : _0315_;
  assign _0317_ = curr_state_r[3] ? opA_r[15] : _0316_;
  assign _0318_ = _0104_ | ~(opA_r[15]);
  assign _0319_ = ~(_0318_ ^ _0317_);
  assign _0320_ = _0302_ | _0301_;
  assign _0321_ = ~(_0309_ | _0303_);
  assign _0322_ = _0320_ & ~(_0321_);
  assign _0323_ = _0322_ ^ _0319_;
  assign _0324_ = gets_high_part_r ? _0323_ : _0310_;
  assign _0325_ = _0040_ ? _0324_ : result_r[15];
  assign _0326_ = ~result_r[14];
  assign _0327_ = _0120_ ? _0326_ : _0310_;
  assign _0717_ = _0039_ ? _0327_ : _0325_;
  assign _0328_ = ~(result_r[16] ^ curr_state_r[1]);
  assign _0329_ = curr_state_r[2] ? opB_r[16] : _0328_;
  assign _0330_ = curr_state_r[3] ? opA_r[16] : _0329_;
  assign _0331_ = _0104_ | ~(opA_r[16]);
  assign _0332_ = ~(_0331_ ^ _0330_);
  assign _0333_ = ~(_0318_ | _0317_);
  assign _0334_ = ~(_0320_ | _0319_);
  assign _0335_ = _0334_ | _0333_;
  assign _0336_ = _0319_ | _0303_;
  assign _0337_ = _0306_ & ~(_0336_);
  assign _0338_ = _0337_ | _0335_;
  assign _0339_ = _0336_ | _0307_;
  assign _0340_ = _0277_ & ~(_0339_);
  assign _0341_ = _0340_ | _0338_;
  assign _0342_ = _0339_ | _0278_;
  assign _0343_ = _0219_ & ~(_0342_);
  assign _0344_ = _0343_ | _0341_;
  assign _0345_ = ~(_0344_ ^ _0332_);
  assign _0346_ = gets_high_part_r ? _0345_ : _0323_;
  assign _0347_ = _0040_ ? _0346_ : result_r[16];
  assign _0348_ = ~result_r[15];
  assign _0349_ = _0120_ ? _0348_ : _0323_;
  assign _0718_ = _0039_ ? _0349_ : _0347_;
  assign _0350_ = ~opA_r[17];
  assign _0351_ = ~opB_r[17];
  assign _0352_ = result_r[17] ^ curr_state_r[1];
  assign _0353_ = curr_state_r[2] ? _0351_ : _0352_;
  assign _0354_ = curr_state_r[3] ? _0350_ : _0353_;
  assign _0355_ = opA_r[17] & ~(_0104_);
  assign _0356_ = _0355_ ^ _0354_;
  assign _0357_ = _0331_ | _0330_;
  assign _0358_ = _0344_ & ~(_0332_);
  assign _0359_ = _0358_ | ~(_0357_);
  assign _0360_ = _0359_ ^ _0356_;
  assign _0361_ = gets_high_part_r ? _0360_ : _0345_;
  assign _0362_ = _0040_ ? _0361_ : result_r[17];
  assign _0363_ = ~result_r[16];
  assign _0364_ = _0120_ ? _0363_ : _0345_;
  assign _0719_ = _0039_ ? _0364_ : _0362_;
  assign _0365_ = ~(result_r[18] ^ curr_state_r[1]);
  assign _0366_ = curr_state_r[2] ? opB_r[18] : _0365_;
  assign _0367_ = curr_state_r[3] ? opA_r[18] : _0366_;
  assign _0368_ = _0104_ | ~(opA_r[18]);
  assign _0369_ = ~(_0368_ ^ _0367_);
  assign _0370_ = _0355_ & _0354_;
  assign _0371_ = _0356_ & ~(_0357_);
  assign _0372_ = _0371_ | _0370_;
  assign _0373_ = _0332_ | ~(_0356_);
  assign _0374_ = _0373_ | ~(_0344_);
  assign _0375_ = _0374_ & ~(_0372_);
  assign _0376_ = _0375_ ^ _0369_;
  assign _0377_ = gets_high_part_r ? _0376_ : _0360_;
  assign _0378_ = _0040_ ? _0377_ : result_r[18];
  assign _0379_ = ~result_r[17];
  assign _0380_ = _0120_ ? _0379_ : _0360_;
  assign _0720_ = _0039_ ? _0380_ : _0378_;
  assign _0381_ = ~(result_r[19] ^ curr_state_r[1]);
  assign _0382_ = curr_state_r[2] ? opB_r[19] : _0381_;
  assign _0383_ = curr_state_r[3] ? opA_r[19] : _0382_;
  assign _0384_ = opA_r[19] & ~(_0104_);
  assign _0385_ = _0384_ ^ _0383_;
  assign _0386_ = _0368_ | _0367_;
  assign _0387_ = ~(_0375_ | _0369_);
  assign _0388_ = _0386_ & ~(_0387_);
  assign _0389_ = _0388_ ^ _0385_;
  assign _0390_ = gets_high_part_r ? _0389_ : _0376_;
  assign _0391_ = _0040_ ? _0390_ : result_r[19];
  assign _0392_ = ~result_r[18];
  assign _0393_ = _0120_ ? _0392_ : _0376_;
  assign _0721_ = _0039_ ? _0393_ : _0391_;
  assign _0394_ = ~(result_r[20] ^ curr_state_r[1]);
  assign _0395_ = curr_state_r[2] ? opB_r[20] : _0394_;
  assign _0396_ = curr_state_r[3] ? opA_r[20] : _0395_;
  assign _0397_ = _0104_ | ~(opA_r[20]);
  assign _0398_ = ~(_0397_ ^ _0396_);
  assign _0399_ = _0384_ & ~(_0383_);
  assign _0400_ = ~(_0386_ | _0385_);
  assign _0401_ = _0400_ | _0399_;
  assign _0402_ = _0385_ | _0369_;
  assign _0403_ = _0372_ & ~(_0402_);
  assign _0404_ = _0403_ | _0401_;
  assign _0405_ = _0402_ | _0373_;
  assign _0406_ = _0344_ & ~(_0405_);
  assign _0407_ = ~(_0406_ | _0404_);
  assign _0408_ = _0407_ ^ _0398_;
  assign _0409_ = gets_high_part_r ? _0408_ : _0389_;
  assign _0410_ = _0040_ ? _0409_ : result_r[20];
  assign _0411_ = ~result_r[19];
  assign _0412_ = _0120_ ? _0411_ : _0389_;
  assign _0722_ = _0039_ ? _0412_ : _0410_;
  assign _0413_ = ~opA_r[21];
  assign _0414_ = ~opB_r[21];
  assign _0415_ = result_r[21] ^ curr_state_r[1];
  assign _0416_ = curr_state_r[2] ? _0414_ : _0415_;
  assign _0417_ = curr_state_r[3] ? _0413_ : _0416_;
  assign _0418_ = opA_r[21] & ~(_0104_);
  assign _0419_ = _0418_ ^ _0417_;
  assign _0420_ = _0397_ | _0396_;
  assign _0421_ = ~(_0407_ | _0398_);
  assign _0422_ = _0421_ | ~(_0420_);
  assign _0423_ = _0422_ ^ _0419_;
  assign _0424_ = gets_high_part_r ? _0423_ : _0408_;
  assign _0425_ = _0040_ ? _0424_ : result_r[21];
  assign _0426_ = ~result_r[20];
  assign _0427_ = _0120_ ? _0426_ : _0408_;
  assign _0724_ = _0039_ ? _0427_ : _0425_;
  assign _0428_ = ~(result_r[22] ^ curr_state_r[1]);
  assign _0429_ = curr_state_r[2] ? opB_r[22] : _0428_;
  assign _0430_ = curr_state_r[3] ? opA_r[22] : _0429_;
  assign _0431_ = opA_r[22] & ~(_0104_);
  assign _0432_ = _0431_ ^ _0430_;
  assign _0433_ = _0418_ & _0417_;
  assign _0434_ = _0419_ & ~(_0420_);
  assign _0435_ = _0434_ | _0433_;
  assign _0436_ = _0398_ | ~(_0419_);
  assign _0437_ = _0436_ | _0407_;
  assign _0438_ = _0437_ & ~(_0435_);
  assign _0439_ = _0438_ ^ _0432_;
  assign _0440_ = gets_high_part_r ? _0439_ : _0423_;
  assign _0441_ = _0040_ ? _0440_ : result_r[22];
  assign _0442_ = ~result_r[21];
  assign _0443_ = _0120_ ? _0442_ : _0423_;
  assign _0725_ = _0039_ ? _0443_ : _0441_;
  assign _0444_ = ~(result_r[23] ^ curr_state_r[1]);
  assign _0445_ = curr_state_r[2] ? opB_r[23] : _0444_;
  assign _0446_ = curr_state_r[3] ? opA_r[23] : _0445_;
  assign _0447_ = opA_r[23] & ~(_0104_);
  assign _0448_ = _0447_ ^ _0446_;
  assign _0449_ = _0430_ | ~(_0431_);
  assign _0450_ = ~(_0438_ | _0432_);
  assign _0451_ = _0449_ & ~(_0450_);
  assign _0452_ = _0451_ ^ _0448_;
  assign _0453_ = gets_high_part_r ? _0452_ : _0439_;
  assign _0454_ = _0040_ ? _0453_ : result_r[23];
  assign _0455_ = ~result_r[22];
  assign _0456_ = _0120_ ? _0455_ : _0439_;
  assign _0726_ = _0039_ ? _0456_ : _0454_;
  assign _0457_ = ~(result_r[24] ^ curr_state_r[1]);
  assign _0458_ = curr_state_r[2] ? opB_r[24] : _0457_;
  assign _0459_ = curr_state_r[3] ? opA_r[24] : _0458_;
  assign _0460_ = opA_r[24] & ~(_0104_);
  assign _0461_ = _0460_ ^ _0459_;
  assign _0462_ = _0447_ & ~(_0446_);
  assign _0463_ = ~(_0449_ | _0448_);
  assign _0464_ = _0463_ | _0462_;
  assign _0465_ = _0448_ | _0432_;
  assign _0466_ = _0435_ & ~(_0465_);
  assign _0467_ = _0466_ | _0464_;
  assign _0468_ = _0465_ | _0436_;
  assign _0469_ = _0404_ & ~(_0468_);
  assign _0470_ = _0469_ | _0467_;
  assign _0471_ = _0468_ | _0405_;
  assign _0472_ = _0344_ & ~(_0471_);
  assign _0473_ = _0472_ | _0470_;
  assign _0474_ = ~(_0473_ ^ _0461_);
  assign _0475_ = gets_high_part_r ? _0474_ : _0452_;
  assign _0476_ = _0040_ ? _0475_ : result_r[24];
  assign _0477_ = ~result_r[23];
  assign _0478_ = _0120_ ? _0477_ : _0452_;
  assign _0727_ = _0039_ ? _0478_ : _0476_;
  assign _0479_ = ~(result_r[25] ^ curr_state_r[1]);
  assign _0480_ = curr_state_r[2] ? opB_r[25] : _0479_;
  assign _0481_ = curr_state_r[3] ? opA_r[25] : _0480_;
  assign _0482_ = opA_r[25] & ~(_0104_);
  assign _0483_ = _0482_ ^ _0481_;
  assign _0484_ = _0459_ | ~(_0460_);
  assign _0485_ = _0473_ & ~(_0461_);
  assign _0486_ = _0484_ & ~(_0485_);
  assign _0487_ = _0486_ ^ _0483_;
  assign _0488_ = gets_high_part_r ? _0487_ : _0474_;
  assign _0489_ = _0040_ ? _0488_ : result_r[25];
  assign _0490_ = ~result_r[24];
  assign _0491_ = _0120_ ? _0490_ : _0474_;
  assign _0728_ = _0039_ ? _0491_ : _0489_;
  assign _0492_ = ~(result_r[26] ^ curr_state_r[1]);
  assign _0493_ = curr_state_r[2] ? opB_r[26] : _0492_;
  assign _0494_ = curr_state_r[3] ? opA_r[26] : _0493_;
  assign _0495_ = opA_r[26] & ~(_0104_);
  assign _0496_ = _0495_ ^ _0494_;
  assign _0497_ = _0482_ & ~(_0481_);
  assign _0498_ = ~(_0484_ | _0483_);
  assign _0499_ = ~(_0498_ | _0497_);
  assign _0500_ = _0483_ | _0461_;
  assign _0501_ = _0473_ & ~(_0500_);
  assign _0502_ = _0499_ & ~(_0501_);
  assign _0503_ = _0502_ ^ _0496_;
  assign _0504_ = gets_high_part_r ? _0503_ : _0487_;
  assign _0505_ = _0040_ ? _0504_ : result_r[26];
  assign _0506_ = ~result_r[25];
  assign _0507_ = _0120_ ? _0506_ : _0487_;
  assign _0729_ = _0039_ ? _0507_ : _0505_;
  assign _0508_ = ~(result_r[27] ^ curr_state_r[1]);
  assign _0509_ = curr_state_r[2] ? opB_r[27] : _0508_;
  assign _0510_ = curr_state_r[3] ? opA_r[27] : _0509_;
  assign _0511_ = opA_r[27] & ~(_0104_);
  assign _0512_ = _0511_ ^ _0510_;
  assign _0513_ = _0494_ | ~(_0495_);
  assign _0514_ = ~(_0502_ | _0496_);
  assign _0515_ = _0513_ & ~(_0514_);
  assign _0516_ = _0515_ ^ _0512_;
  assign _0517_ = gets_high_part_r ? _0516_ : _0503_;
  assign _0518_ = _0040_ ? _0517_ : result_r[27];
  assign _0519_ = ~result_r[26];
  assign _0520_ = _0120_ ? _0519_ : _0503_;
  assign _0730_ = _0039_ ? _0520_ : _0518_;
  assign _0521_ = ~(result_r[28] ^ curr_state_r[1]);
  assign _0522_ = curr_state_r[2] ? opB_r[28] : _0521_;
  assign _0523_ = curr_state_r[3] ? opA_r[28] : _0522_;
  assign _0524_ = opA_r[28] & ~(_0104_);
  assign _0525_ = _0524_ ^ _0523_;
  assign _0526_ = _0511_ & ~(_0510_);
  assign _0527_ = ~(_0513_ | _0512_);
  assign _0528_ = _0527_ | _0526_;
  assign _0529_ = _0512_ | _0496_;
  assign _0530_ = ~(_0529_ | _0499_);
  assign _0531_ = _0530_ | _0528_;
  assign _0532_ = _0529_ | _0500_;
  assign _0533_ = _0473_ & ~(_0532_);
  assign _0534_ = ~(_0533_ | _0531_);
  assign _0535_ = _0534_ ^ _0525_;
  assign _0536_ = gets_high_part_r ? _0535_ : _0516_;
  assign _0537_ = _0040_ ? _0536_ : result_r[28];
  assign _0538_ = ~result_r[27];
  assign _0539_ = _0120_ ? _0538_ : _0516_;
  assign _0731_ = _0039_ ? _0539_ : _0537_;
  assign _0540_ = ~(result_r[29] ^ curr_state_r[1]);
  assign _0541_ = curr_state_r[2] ? opB_r[29] : _0540_;
  assign _0542_ = curr_state_r[3] ? opA_r[29] : _0541_;
  assign _0543_ = opA_r[29] & ~(_0104_);
  assign _0544_ = _0543_ ^ _0542_;
  assign _0545_ = _0523_ | ~(_0524_);
  assign _0546_ = ~(_0534_ | _0525_);
  assign _0547_ = _0545_ & ~(_0546_);
  assign _0548_ = _0547_ ^ _0544_;
  assign _0549_ = gets_high_part_r ? _0548_ : _0535_;
  assign _0550_ = _0040_ ? _0549_ : result_r[29];
  assign _0551_ = ~result_r[28];
  assign _0552_ = _0120_ ? _0551_ : _0535_;
  assign _0732_ = _0039_ ? _0552_ : _0550_;
  assign _0553_ = ~(result_r[30] ^ curr_state_r[1]);
  assign _0554_ = curr_state_r[2] ? opB_r[30] : _0553_;
  assign _0555_ = curr_state_r[3] ? opA_r[30] : _0554_;
  assign _0556_ = opA_r[30] & ~(_0104_);
  assign _0557_ = _0556_ ^ _0555_;
  assign _0558_ = _0543_ & ~(_0542_);
  assign _0559_ = ~(_0545_ | _0544_);
  assign _0560_ = ~(_0559_ | _0558_);
  assign _0561_ = _0544_ | _0525_;
  assign _0562_ = ~(_0561_ | _0534_);
  assign _0563_ = _0560_ & ~(_0562_);
  assign _0564_ = _0563_ ^ _0557_;
  assign _0565_ = gets_high_part_r ? _0564_ : _0548_;
  assign _0566_ = _0040_ ? _0565_ : result_r[30];
  assign _0567_ = ~result_r[29];
  assign _0568_ = _0120_ ? _0567_ : _0548_;
  assign _0733_ = _0039_ ? _0568_ : _0566_;
  assign _0569_ = ~(result_r[31] ^ curr_state_r[1]);
  assign _0570_ = curr_state_r[2] ? opB_r[31] : _0569_;
  assign _0571_ = curr_state_r[3] ? opA_r[31] : _0570_;
  assign _0572_ = opA_r[31] & ~(_0104_);
  assign _0573_ = _0572_ ^ _0571_;
  assign _0574_ = _0555_ | ~(_0556_);
  assign _0575_ = ~(_0563_ | _0557_);
  assign _0576_ = _0574_ & ~(_0575_);
  assign _0577_ = _0576_ ^ _0573_;
  assign _0578_ = gets_high_part_r ? _0577_ : _0564_;
  assign _0579_ = _0040_ ? _0578_ : result_r[31];
  assign _0580_ = ~result_r[30];
  assign _0581_ = _0120_ ? _0580_ : _0564_;
  assign _0735_ = _0039_ ? _0581_ : _0579_;
  assign _0582_ = ~(_0576_ ^ _0573_);
  assign _0583_ = _0571_ | ~(_0572_);
  assign _0584_ = ~(_0574_ | _0573_);
  assign _0585_ = _0583_ & ~(_0584_);
  assign _0586_ = _0573_ | _0557_;
  assign _0587_ = ~(_0586_ | _0560_);
  assign _0588_ = _0585_ & ~(_0587_);
  assign _0589_ = _0586_ | _0561_;
  assign _0590_ = _0531_ & ~(_0589_);
  assign _0591_ = _0588_ & ~(_0590_);
  assign _0592_ = _0589_ | _0532_;
  assign _0593_ = _0470_ & ~(_0592_);
  assign _0594_ = _0591_ & ~(_0593_);
  assign _0595_ = _0592_ | _0471_;
  assign _0596_ = _0344_ & ~(_0595_);
  assign _0597_ = _0594_ & ~(_0596_);
  assign _0598_ = gets_high_part_r ? _0597_ : _0582_;
  assign _0599_ = ~(_0598_ | _0100_);
  assign _0600_ = ~result_r[31];
  assign _0601_ = _0120_ ? _0600_ : _0577_;
  assign _0736_ = _0039_ ? _0601_ : _0599_;
  assign _0602_ = curr_state_r[5] ? opB_r[1] : _0107_;
  assign _0648_ = latch_input ? opB_i[0] : _0602_;
  assign _0603_ = curr_state_r[5] ? opB_r[2] : _0116_;
  assign _0659_ = latch_input ? opB_i[1] : _0603_;
  assign _0604_ = curr_state_r[5] ? opB_r[3] : _0130_;
  assign _0670_ = latch_input ? opB_i[2] : _0604_;
  assign _0605_ = curr_state_r[5] ? opB_r[4] : _0143_;
  assign _0673_ = latch_input ? opB_i[3] : _0605_;
  assign _0606_ = curr_state_r[5] ? opB_r[5] : _0159_;
  assign _0674_ = latch_input ? opB_i[4] : _0606_;
  assign _0607_ = curr_state_r[5] ? opB_r[6] : _0172_;
  assign _0675_ = latch_input ? opB_i[5] : _0607_;
  assign _0608_ = curr_state_r[5] ? opB_r[7] : _0188_;
  assign _0676_ = latch_input ? opB_i[6] : _0608_;
  assign _0609_ = curr_state_r[5] ? opB_r[8] : _0201_;
  assign _0677_ = latch_input ? opB_i[7] : _0609_;
  assign _0610_ = curr_state_r[5] ? opB_r[9] : _0220_;
  assign _0678_ = latch_input ? opB_i[8] : _0610_;
  assign _0611_ = curr_state_r[5] ? opB_r[10] : _0233_;
  assign _0679_ = latch_input ? opB_i[9] : _0611_;
  assign _0612_ = curr_state_r[5] ? opB_r[11] : _0249_;
  assign _0649_ = latch_input ? opB_i[10] : _0612_;
  assign _0613_ = curr_state_r[5] ? opB_r[12] : _0262_;
  assign _0650_ = latch_input ? opB_i[11] : _0613_;
  assign _0614_ = curr_state_r[5] ? opB_r[13] : _0281_;
  assign _0651_ = latch_input ? opB_i[12] : _0614_;
  assign _0615_ = curr_state_r[5] ? opB_r[14] : _0294_;
  assign _0652_ = latch_input ? opB_i[13] : _0615_;
  assign _0616_ = curr_state_r[5] ? opB_r[15] : _0310_;
  assign _0653_ = latch_input ? opB_i[14] : _0616_;
  assign _0617_ = curr_state_r[5] ? opB_r[16] : _0323_;
  assign _0654_ = latch_input ? opB_i[15] : _0617_;
  assign _0618_ = curr_state_r[5] ? opB_r[17] : _0345_;
  assign _0655_ = latch_input ? opB_i[16] : _0618_;
  assign _0619_ = curr_state_r[5] ? opB_r[18] : _0360_;
  assign _0656_ = latch_input ? opB_i[17] : _0619_;
  assign _0620_ = curr_state_r[5] ? opB_r[19] : _0376_;
  assign _0657_ = latch_input ? opB_i[18] : _0620_;
  assign _0621_ = curr_state_r[5] ? opB_r[20] : _0389_;
  assign _0658_ = latch_input ? opB_i[19] : _0621_;
  assign _0622_ = curr_state_r[5] ? opB_r[21] : _0408_;
  assign _0660_ = latch_input ? opB_i[20] : _0622_;
  assign _0623_ = curr_state_r[5] ? opB_r[22] : _0423_;
  assign _0661_ = latch_input ? opB_i[21] : _0623_;
  assign _0624_ = curr_state_r[5] ? opB_r[23] : _0439_;
  assign _0662_ = latch_input ? opB_i[22] : _0624_;
  assign _0625_ = curr_state_r[5] ? opB_r[24] : _0452_;
  assign _0663_ = latch_input ? opB_i[23] : _0625_;
  assign _0626_ = curr_state_r[5] ? opB_r[25] : _0474_;
  assign _0664_ = latch_input ? opB_i[24] : _0626_;
  assign _0627_ = curr_state_r[5] ? opB_r[26] : _0487_;
  assign _0665_ = latch_input ? opB_i[25] : _0627_;
  assign _0628_ = curr_state_r[5] ? opB_r[27] : _0503_;
  assign _0666_ = latch_input ? opB_i[26] : _0628_;
  assign _0629_ = curr_state_r[5] ? opB_r[28] : _0516_;
  assign _0667_ = latch_input ? opB_i[27] : _0629_;
  assign _0630_ = curr_state_r[5] ? opB_r[29] : _0535_;
  assign _0668_ = latch_input ? opB_i[28] : _0630_;
  assign _0631_ = curr_state_r[5] ? opB_r[30] : _0548_;
  assign _0669_ = latch_input ? opB_i[29] : _0631_;
  assign _0632_ = curr_state_r[5] ? opB_r[31] : _0564_;
  assign _0671_ = latch_input ? opB_i[30] : _0632_;
  assign _0633_ = _0086_ & ~(_0582_);
  assign _0672_ = latch_input ? opB_i[31] : _0633_;
  assign _0634_ = ~(_0106_ | _0097_);
  assign _0680_ = latch_input ? opA_i[0] : _0634_;
  assign _0635_ = _0097_ ? opA_r[0] : _0116_;
  assign _0691_ = latch_input ? opA_i[1] : _0635_;
  assign _0636_ = _0097_ ? opA_r[1] : _0130_;
  assign _0702_ = latch_input ? opA_i[2] : _0636_;
  assign _0637_ = _0097_ ? opA_r[2] : _0143_;
  assign _0705_ = latch_input ? opA_i[3] : _0637_;
  assign _0638_ = _0097_ ? opA_r[3] : _0159_;
  assign _0706_ = latch_input ? opA_i[4] : _0638_;
  assign _0639_ = _0097_ ? opA_r[4] : _0172_;
  assign _0707_ = latch_input ? opA_i[5] : _0639_;
  assign _0640_ = _0097_ ? opA_r[5] : _0188_;
  assign _0708_ = latch_input ? opA_i[6] : _0640_;
  assign _0641_ = _0097_ ? opA_r[6] : _0201_;
  assign _0709_ = latch_input ? opA_i[7] : _0641_;
  assign _0642_ = _0097_ ? opA_r[7] : _0220_;
  assign _0710_ = latch_input ? opA_i[8] : _0642_;
  assign _0643_ = _0097_ ? opA_r[8] : _0233_;
  assign _0711_ = latch_input ? opA_i[9] : _0643_;
  assign _0644_ = _0097_ ? opA_r[9] : _0249_;
  assign _0681_ = latch_input ? opA_i[10] : _0644_;
  assign _0645_ = _0097_ ? opA_r[10] : _0262_;
  assign _0682_ = latch_input ? opA_i[11] : _0645_;
  assign _0646_ = _0097_ ? opA_r[11] : _0281_;
  assign _0683_ = latch_input ? opA_i[12] : _0646_;
  assign _0647_ = _0097_ ? opA_r[12] : _0294_;
  assign _0684_ = latch_input ? opA_i[13] : _0647_;
  assign _0012_ = _0097_ ? opA_r[13] : _0310_;
  assign _0685_ = latch_input ? opA_i[14] : _0012_;
  assign _0013_ = _0097_ ? opA_r[14] : _0323_;
  assign _0686_ = latch_input ? opA_i[15] : _0013_;
  assign _0014_ = _0097_ ? opA_r[15] : _0345_;
  assign _0687_ = latch_input ? opA_i[16] : _0014_;
  assign _0015_ = _0097_ ? opA_r[16] : _0360_;
  assign _0688_ = latch_input ? opA_i[17] : _0015_;
  assign _0016_ = _0097_ ? opA_r[17] : _0376_;
  assign _0689_ = latch_input ? opA_i[18] : _0016_;
  assign _0017_ = _0097_ ? opA_r[18] : _0389_;
  assign _0690_ = latch_input ? opA_i[19] : _0017_;
  assign _0018_ = _0097_ ? opA_r[19] : _0408_;
  assign _0692_ = latch_input ? opA_i[20] : _0018_;
  assign _0019_ = _0097_ ? opA_r[20] : _0423_;
  assign _0693_ = latch_input ? opA_i[21] : _0019_;
  assign _0020_ = _0097_ ? opA_r[21] : _0439_;
  assign _0694_ = latch_input ? opA_i[22] : _0020_;
  assign _0021_ = _0097_ ? opA_r[22] : _0452_;
  assign _0695_ = latch_input ? opA_i[23] : _0021_;
  assign _0022_ = _0097_ ? opA_r[23] : _0474_;
  assign _0696_ = latch_input ? opA_i[24] : _0022_;
  assign _0023_ = _0097_ ? opA_r[24] : _0487_;
  assign _0697_ = latch_input ? opA_i[25] : _0023_;
  assign _0024_ = _0097_ ? opA_r[25] : _0503_;
  assign _0698_ = latch_input ? opA_i[26] : _0024_;
  assign _0025_ = _0097_ ? opA_r[26] : _0516_;
  assign _0699_ = latch_input ? opA_i[27] : _0025_;
  assign _0026_ = _0097_ ? opA_r[27] : _0535_;
  assign _0700_ = latch_input ? opA_i[28] : _0026_;
  assign _0027_ = _0097_ ? opA_r[28] : _0548_;
  assign _0701_ = latch_input ? opA_i[29] : _0027_;
  assign _0028_ = _0097_ ? opA_r[29] : _0564_;
  assign _0703_ = latch_input ? opA_i[30] : _0028_;
  assign _0029_ = _0097_ ? opA_r[30] : _0577_;
  assign _0704_ = latch_input ? opA_i[31] : _0029_;
  assign _0747_[1] = shift_counter_r[1] ^ shift_counter_r[0];
  assign _0030_ = shift_counter_r[1] & shift_counter_r[0];
  assign _0747_[2] = _0030_ ^ shift_counter_r[2];
  assign _0031_ = _0030_ & shift_counter_r[2];
  assign _0747_[3] = _0031_ ^ shift_counter_r[3];
  assign _0032_ = ~(shift_counter_r[3] & shift_counter_r[2]);
  assign _0033_ = _0030_ & ~(_0032_);
  assign _0747_[4] = _0033_ ^ shift_counter_r[4];
  assign _0034_ = _0033_ & shift_counter_r[4];
  assign _0747_[5] = _0034_ ^ shift_counter_r[5];
  assign signed_opA = signed_opA_i & opA_i[31];
  assign signed_opB = signed_opB_i & opB_i[31];
  assign _0745_ = signed_opB ^ signed_opA;
  assign _0035_ = reset_i | ~(_0072_);
  assign _0000_ = curr_state_r[5] & ~(_0035_);
  assign _0036_ = opB_r[0] ? _0106_ : _0119_;
  assign _0037_ = _0036_ & all_sh_lsb_zero_r;
  assign _0744_ = _0037_ | latch_input;
  assign _0001_ = curr_state_r[3] & ~(reset_i);
  assign _0038_ = reset_i | ~(v_i);
  assign _0002_ = curr_state_r[0] & ~(_0038_);
  always @(posedge clk_i)
    if (_0009_) result_r[0] <= 1'h0;
    else if (_0007_) result_r[0] <= _0712_;
  always @(posedge clk_i)
    if (_0009_) result_r[1] <= 1'h0;
    else if (_0007_) result_r[1] <= _0723_;
  always @(posedge clk_i)
    if (_0009_) result_r[2] <= 1'h0;
    else if (_0007_) result_r[2] <= _0734_;
  always @(posedge clk_i)
    if (_0009_) result_r[3] <= 1'h0;
    else if (_0007_) result_r[3] <= _0737_;
  always @(posedge clk_i)
    if (_0009_) result_r[4] <= 1'h0;
    else if (_0007_) result_r[4] <= _0738_;
  always @(posedge clk_i)
    if (_0009_) result_r[5] <= 1'h0;
    else if (_0007_) result_r[5] <= _0739_;
  always @(posedge clk_i)
    if (_0009_) result_r[6] <= 1'h0;
    else if (_0007_) result_r[6] <= _0740_;
  always @(posedge clk_i)
    if (_0009_) result_r[7] <= 1'h0;
    else if (_0007_) result_r[7] <= _0741_;
  always @(posedge clk_i)
    if (_0009_) result_r[8] <= 1'h0;
    else if (_0007_) result_r[8] <= _0742_;
  always @(posedge clk_i)
    if (_0009_) result_r[9] <= 1'h0;
    else if (_0007_) result_r[9] <= _0743_;
  always @(posedge clk_i)
    if (_0009_) result_r[10] <= 1'h0;
    else if (_0007_) result_r[10] <= _0713_;
  always @(posedge clk_i)
    if (_0009_) result_r[11] <= 1'h0;
    else if (_0007_) result_r[11] <= _0714_;
  always @(posedge clk_i)
    if (_0009_) result_r[12] <= 1'h0;
    else if (_0007_) result_r[12] <= _0715_;
  always @(posedge clk_i)
    if (_0009_) result_r[13] <= 1'h0;
    else if (_0007_) result_r[13] <= _0716_;
  always @(posedge clk_i)
    if (_0009_) result_r[14] <= 1'h0;
    else if (_0007_) result_r[14] <= _0717_;
  always @(posedge clk_i)
    if (_0009_) result_r[15] <= 1'h0;
    else if (_0007_) result_r[15] <= _0718_;
  always @(posedge clk_i)
    if (_0009_) result_r[16] <= 1'h0;
    else if (_0007_) result_r[16] <= _0719_;
  always @(posedge clk_i)
    if (_0009_) result_r[17] <= 1'h0;
    else if (_0007_) result_r[17] <= _0720_;
  always @(posedge clk_i)
    if (_0009_) result_r[18] <= 1'h0;
    else if (_0007_) result_r[18] <= _0721_;
  always @(posedge clk_i)
    if (_0009_) result_r[19] <= 1'h0;
    else if (_0007_) result_r[19] <= _0722_;
  always @(posedge clk_i)
    if (_0009_) result_r[20] <= 1'h0;
    else if (_0007_) result_r[20] <= _0724_;
  always @(posedge clk_i)
    if (_0009_) result_r[21] <= 1'h0;
    else if (_0007_) result_r[21] <= _0725_;
  always @(posedge clk_i)
    if (_0009_) result_r[22] <= 1'h0;
    else if (_0007_) result_r[22] <= _0726_;
  always @(posedge clk_i)
    if (_0009_) result_r[23] <= 1'h0;
    else if (_0007_) result_r[23] <= _0727_;
  always @(posedge clk_i)
    if (_0009_) result_r[24] <= 1'h0;
    else if (_0007_) result_r[24] <= _0728_;
  always @(posedge clk_i)
    if (_0009_) result_r[25] <= 1'h0;
    else if (_0007_) result_r[25] <= _0729_;
  always @(posedge clk_i)
    if (_0009_) result_r[26] <= 1'h0;
    else if (_0007_) result_r[26] <= _0730_;
  always @(posedge clk_i)
    if (_0009_) result_r[27] <= 1'h0;
    else if (_0007_) result_r[27] <= _0731_;
  always @(posedge clk_i)
    if (_0009_) result_r[28] <= 1'h0;
    else if (_0007_) result_r[28] <= _0732_;
  always @(posedge clk_i)
    if (_0009_) result_r[29] <= 1'h0;
    else if (_0007_) result_r[29] <= _0733_;
  always @(posedge clk_i)
    if (_0009_) result_r[30] <= 1'h0;
    else if (_0007_) result_r[30] <= _0735_;
  always @(posedge clk_i)
    if (_0009_) result_r[31] <= 1'h0;
    else if (_0007_) result_r[31] <= _0736_;
  always @(posedge clk_i)
    if (reset_i) all_sh_lsb_zero_r <= 1'h0;
    else if (_0006_) all_sh_lsb_zero_r <= _0744_;
  always @(posedge clk_i)
    if (reset_i) opB_r[0] <= 1'h0;
    else if (_0005_) opB_r[0] <= _0648_;
  always @(posedge clk_i)
    if (reset_i) opB_r[1] <= 1'h0;
    else if (_0005_) opB_r[1] <= _0659_;
  always @(posedge clk_i)
    if (reset_i) opB_r[2] <= 1'h0;
    else if (_0005_) opB_r[2] <= _0670_;
  always @(posedge clk_i)
    if (reset_i) opB_r[3] <= 1'h0;
    else if (_0005_) opB_r[3] <= _0673_;
  always @(posedge clk_i)
    if (reset_i) opB_r[4] <= 1'h0;
    else if (_0005_) opB_r[4] <= _0674_;
  always @(posedge clk_i)
    if (reset_i) opB_r[5] <= 1'h0;
    else if (_0005_) opB_r[5] <= _0675_;
  always @(posedge clk_i)
    if (reset_i) opB_r[6] <= 1'h0;
    else if (_0005_) opB_r[6] <= _0676_;
  always @(posedge clk_i)
    if (reset_i) opB_r[7] <= 1'h0;
    else if (_0005_) opB_r[7] <= _0677_;
  always @(posedge clk_i)
    if (reset_i) opB_r[8] <= 1'h0;
    else if (_0005_) opB_r[8] <= _0678_;
  always @(posedge clk_i)
    if (reset_i) opB_r[9] <= 1'h0;
    else if (_0005_) opB_r[9] <= _0679_;
  always @(posedge clk_i)
    if (reset_i) opB_r[10] <= 1'h0;
    else if (_0005_) opB_r[10] <= _0649_;
  always @(posedge clk_i)
    if (reset_i) opB_r[11] <= 1'h0;
    else if (_0005_) opB_r[11] <= _0650_;
  always @(posedge clk_i)
    if (reset_i) opB_r[12] <= 1'h0;
    else if (_0005_) opB_r[12] <= _0651_;
  always @(posedge clk_i)
    if (reset_i) opB_r[13] <= 1'h0;
    else if (_0005_) opB_r[13] <= _0652_;
  always @(posedge clk_i)
    if (reset_i) opB_r[14] <= 1'h0;
    else if (_0005_) opB_r[14] <= _0653_;
  always @(posedge clk_i)
    if (reset_i) opB_r[15] <= 1'h0;
    else if (_0005_) opB_r[15] <= _0654_;
  always @(posedge clk_i)
    if (reset_i) opB_r[16] <= 1'h0;
    else if (_0005_) opB_r[16] <= _0655_;
  always @(posedge clk_i)
    if (reset_i) opB_r[17] <= 1'h0;
    else if (_0005_) opB_r[17] <= _0656_;
  always @(posedge clk_i)
    if (reset_i) opB_r[18] <= 1'h0;
    else if (_0005_) opB_r[18] <= _0657_;
  always @(posedge clk_i)
    if (reset_i) opB_r[19] <= 1'h0;
    else if (_0005_) opB_r[19] <= _0658_;
  always @(posedge clk_i)
    if (reset_i) opB_r[20] <= 1'h0;
    else if (_0005_) opB_r[20] <= _0660_;
  always @(posedge clk_i)
    if (reset_i) opB_r[21] <= 1'h0;
    else if (_0005_) opB_r[21] <= _0661_;
  always @(posedge clk_i)
    if (reset_i) opB_r[22] <= 1'h0;
    else if (_0005_) opB_r[22] <= _0662_;
  always @(posedge clk_i)
    if (reset_i) opB_r[23] <= 1'h0;
    else if (_0005_) opB_r[23] <= _0663_;
  always @(posedge clk_i)
    if (reset_i) opB_r[24] <= 1'h0;
    else if (_0005_) opB_r[24] <= _0664_;
  always @(posedge clk_i)
    if (reset_i) opB_r[25] <= 1'h0;
    else if (_0005_) opB_r[25] <= _0665_;
  always @(posedge clk_i)
    if (reset_i) opB_r[26] <= 1'h0;
    else if (_0005_) opB_r[26] <= _0666_;
  always @(posedge clk_i)
    if (reset_i) opB_r[27] <= 1'h0;
    else if (_0005_) opB_r[27] <= _0667_;
  always @(posedge clk_i)
    if (reset_i) opB_r[28] <= 1'h0;
    else if (_0005_) opB_r[28] <= _0668_;
  always @(posedge clk_i)
    if (reset_i) opB_r[29] <= 1'h0;
    else if (_0005_) opB_r[29] <= _0669_;
  always @(posedge clk_i)
    if (reset_i) opB_r[30] <= 1'h0;
    else if (_0005_) opB_r[30] <= _0671_;
  always @(posedge clk_i)
    if (reset_i) opB_r[31] <= 1'h0;
    else if (_0005_) opB_r[31] <= _0672_;
  always @(posedge clk_i)
    if (reset_i) opA_r[0] <= 1'h0;
    else if (_0004_) opA_r[0] <= _0680_;
  always @(posedge clk_i)
    if (reset_i) opA_r[1] <= 1'h0;
    else if (_0004_) opA_r[1] <= _0691_;
  always @(posedge clk_i)
    if (reset_i) opA_r[2] <= 1'h0;
    else if (_0004_) opA_r[2] <= _0702_;
  always @(posedge clk_i)
    if (reset_i) opA_r[3] <= 1'h0;
    else if (_0004_) opA_r[3] <= _0705_;
  always @(posedge clk_i)
    if (reset_i) opA_r[4] <= 1'h0;
    else if (_0004_) opA_r[4] <= _0706_;
  always @(posedge clk_i)
    if (reset_i) opA_r[5] <= 1'h0;
    else if (_0004_) opA_r[5] <= _0707_;
  always @(posedge clk_i)
    if (reset_i) opA_r[6] <= 1'h0;
    else if (_0004_) opA_r[6] <= _0708_;
  always @(posedge clk_i)
    if (reset_i) opA_r[7] <= 1'h0;
    else if (_0004_) opA_r[7] <= _0709_;
  always @(posedge clk_i)
    if (reset_i) opA_r[8] <= 1'h0;
    else if (_0004_) opA_r[8] <= _0710_;
  always @(posedge clk_i)
    if (reset_i) opA_r[9] <= 1'h0;
    else if (_0004_) opA_r[9] <= _0711_;
  always @(posedge clk_i)
    if (reset_i) opA_r[10] <= 1'h0;
    else if (_0004_) opA_r[10] <= _0681_;
  always @(posedge clk_i)
    if (reset_i) opA_r[11] <= 1'h0;
    else if (_0004_) opA_r[11] <= _0682_;
  always @(posedge clk_i)
    if (reset_i) opA_r[12] <= 1'h0;
    else if (_0004_) opA_r[12] <= _0683_;
  always @(posedge clk_i)
    if (reset_i) opA_r[13] <= 1'h0;
    else if (_0004_) opA_r[13] <= _0684_;
  always @(posedge clk_i)
    if (reset_i) opA_r[14] <= 1'h0;
    else if (_0004_) opA_r[14] <= _0685_;
  always @(posedge clk_i)
    if (reset_i) opA_r[15] <= 1'h0;
    else if (_0004_) opA_r[15] <= _0686_;
  always @(posedge clk_i)
    if (reset_i) opA_r[16] <= 1'h0;
    else if (_0004_) opA_r[16] <= _0687_;
  always @(posedge clk_i)
    if (reset_i) opA_r[17] <= 1'h0;
    else if (_0004_) opA_r[17] <= _0688_;
  always @(posedge clk_i)
    if (reset_i) opA_r[18] <= 1'h0;
    else if (_0004_) opA_r[18] <= _0689_;
  always @(posedge clk_i)
    if (reset_i) opA_r[19] <= 1'h0;
    else if (_0004_) opA_r[19] <= _0690_;
  always @(posedge clk_i)
    if (reset_i) opA_r[20] <= 1'h0;
    else if (_0004_) opA_r[20] <= _0692_;
  always @(posedge clk_i)
    if (reset_i) opA_r[21] <= 1'h0;
    else if (_0004_) opA_r[21] <= _0693_;
  always @(posedge clk_i)
    if (reset_i) opA_r[22] <= 1'h0;
    else if (_0004_) opA_r[22] <= _0694_;
  always @(posedge clk_i)
    if (reset_i) opA_r[23] <= 1'h0;
    else if (_0004_) opA_r[23] <= _0695_;
  always @(posedge clk_i)
    if (reset_i) opA_r[24] <= 1'h0;
    else if (_0004_) opA_r[24] <= _0696_;
  always @(posedge clk_i)
    if (reset_i) opA_r[25] <= 1'h0;
    else if (_0004_) opA_r[25] <= _0697_;
  always @(posedge clk_i)
    if (reset_i) opA_r[26] <= 1'h0;
    else if (_0004_) opA_r[26] <= _0698_;
  always @(posedge clk_i)
    if (reset_i) opA_r[27] <= 1'h0;
    else if (_0004_) opA_r[27] <= _0699_;
  always @(posedge clk_i)
    if (reset_i) opA_r[28] <= 1'h0;
    else if (_0004_) opA_r[28] <= _0700_;
  always @(posedge clk_i)
    if (reset_i) opA_r[29] <= 1'h0;
    else if (_0004_) opA_r[29] <= _0701_;
  always @(posedge clk_i)
    if (reset_i) opA_r[30] <= 1'h0;
    else if (_0004_) opA_r[30] <= _0703_;
  always @(posedge clk_i)
    if (reset_i) opA_r[31] <= 1'h0;
    else if (_0004_) opA_r[31] <= _0704_;
  always @(posedge clk_i)
    if (reset_i) gets_high_part_r <= 1'h0;
    else if (latch_input) gets_high_part_r <= gets_high_part_i;
  always @(posedge clk_i)
    if (reset_i) need_neg_result_r <= 1'h0;
    else if (latch_input) need_neg_result_r <= _0745_;
  always @(posedge clk_i)
    if (reset_i) signed_opB_r <= 1'h0;
    else if (latch_input) signed_opB_r <= signed_opB;
  always @(posedge clk_i)
    if (reset_i) signed_opA_r <= 1'h0;
    else if (latch_input) signed_opA_r <= signed_opA;
  always @(posedge clk_i)
    if (_0008_) shift_counter_r[0] <= 1'h0;
    else if (curr_state_r[5]) shift_counter_r[0] <= _0746_[0];
  always @(posedge clk_i)
    if (_0008_) shift_counter_r[1] <= 1'h0;
    else if (curr_state_r[5]) shift_counter_r[1] <= _0747_[1];
  always @(posedge clk_i)
    if (_0008_) shift_counter_r[2] <= 1'h0;
    else if (curr_state_r[5]) shift_counter_r[2] <= _0747_[2];
  always @(posedge clk_i)
    if (_0008_) shift_counter_r[3] <= 1'h0;
    else if (curr_state_r[5]) shift_counter_r[3] <= _0747_[3];
  always @(posedge clk_i)
    if (_0008_) shift_counter_r[4] <= 1'h0;
    else if (curr_state_r[5]) shift_counter_r[4] <= _0747_[4];
  always @(posedge clk_i)
    if (_0008_) shift_counter_r[5] <= 1'h0;
    else if (curr_state_r[5]) shift_counter_r[5] <= _0747_[5];
  always @(posedge clk_i)
    curr_state_r[0] <= _0003_;
  always @(posedge clk_i)
    curr_state_r[1] <= _0000_;
  always @(posedge clk_i)
    curr_state_r[2] <= _0001_;
  always @(posedge clk_i)
    curr_state_r[3] <= _0002_;
  always @(posedge clk_i)
    curr_state_r[4] <= _0010_;
  always @(posedge clk_i)
    curr_state_r[5] <= _0011_;
  assign _0746_[5:1] = shift_counter_r[5:1];
  assign _0747_[0] = _0746_[0];
  assign ready_o = curr_state_r[0];
  assign result_o = result_r;
  assign v_o = curr_state_r[4];
endmodule
