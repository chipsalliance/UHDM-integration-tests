module bsg_round_robin_1_to_n(clk_i, reset_i, valid_i, ready_o, valid_o, ready_i);
  input clk_i;
  wire clk_i;
  wire \one_to_n.circular_ptr.add_i ;
  wire \one_to_n.circular_ptr.clk ;
  wire \one_to_n.circular_ptr.genblk1.genblk1.ptr_r_p1 ;
  wire \one_to_n.circular_ptr.o ;
  reg \one_to_n.circular_ptr.ptr_r ;
  wire \one_to_n.circular_ptr.reset_i ;
  wire \one_to_n.ptr_r ;
  wire \one_to_n.yumi_i ;
  input [1:0] ready_i;
  wire [1:0] ready_i;
  output ready_o;
  wire ready_o;
  input reset_i;
  wire reset_i;
  input valid_i;
  wire valid_i;
  output [1:0] valid_o;
  wire [1:0] valid_o;
  assign \one_to_n.circular_ptr.genblk1.genblk1.ptr_r_p1  = ~\one_to_n.circular_ptr.ptr_r ;
  assign ready_o = \one_to_n.circular_ptr.ptr_r  ? ready_i[1] : ready_i[0];
  assign \one_to_n.circular_ptr.add_i  = ready_o & valid_i;
  assign valid_o[0] = valid_i & ~(\one_to_n.circular_ptr.ptr_r );
  assign valid_o[1] = valid_i & \one_to_n.circular_ptr.ptr_r ;
  always @(posedge clk_i)
    if (reset_i) \one_to_n.circular_ptr.ptr_r  <= 1'h0;
    else if (\one_to_n.circular_ptr.add_i ) \one_to_n.circular_ptr.ptr_r  <= \one_to_n.circular_ptr.genblk1.genblk1.ptr_r_p1 ;
  assign \one_to_n.circular_ptr.clk  = clk_i;
  assign \one_to_n.circular_ptr.o  = \one_to_n.circular_ptr.ptr_r ;
  assign \one_to_n.circular_ptr.reset_i  = reset_i;
  assign \one_to_n.ptr_r  = \one_to_n.circular_ptr.ptr_r ;
  assign \one_to_n.yumi_i  = \one_to_n.circular_ptr.add_i ;
endmodule
