module bsg_permute_box(data_i, select_i, data_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  input [15:0] data_i;
  wire [15:0] data_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  input [31:0] select_i;
  wire [31:0] select_i;
  assign _00_ = ~select_i[0];
  assign _01_ = select_i[1] | ~(data_i[0]);
  assign data_o[0] = _00_ & ~(_01_);
  assign _02_ = select_i[1] | ~(data_i[1]);
  assign data_o[1] = _00_ & ~(_02_);
  assign _03_ = select_i[1] | ~(data_i[2]);
  assign data_o[2] = _00_ & ~(_03_);
  assign _04_ = select_i[1] | ~(data_i[3]);
  assign data_o[3] = _00_ & ~(_04_);
  assign _05_ = select_i[1] | ~(data_i[4]);
  assign data_o[4] = _00_ & ~(_05_);
  assign _06_ = select_i[1] | ~(data_i[5]);
  assign data_o[5] = _00_ & ~(_06_);
  assign _07_ = select_i[1] | ~(data_i[6]);
  assign data_o[6] = _00_ & ~(_07_);
  assign _08_ = select_i[1] | ~(data_i[7]);
  assign data_o[7] = _00_ & ~(_08_);
  assign _09_ = select_i[1] | ~(data_i[8]);
  assign data_o[8] = _00_ & ~(_09_);
  assign _10_ = select_i[1] | ~(data_i[9]);
  assign data_o[9] = _00_ & ~(_10_);
  assign _11_ = select_i[1] | ~(data_i[10]);
  assign data_o[10] = _00_ & ~(_11_);
  assign _12_ = select_i[1] | ~(data_i[11]);
  assign data_o[11] = _00_ & ~(_12_);
  assign _13_ = select_i[1] | ~(data_i[12]);
  assign data_o[12] = _00_ & ~(_13_);
  assign _14_ = select_i[1] | ~(data_i[13]);
  assign data_o[13] = _00_ & ~(_14_);
  assign _15_ = select_i[1] | ~(data_i[14]);
  assign data_o[14] = _00_ & ~(_15_);
  assign _16_ = select_i[1] | ~(data_i[15]);
  assign data_o[15] = _00_ & ~(_16_);
endmodule
