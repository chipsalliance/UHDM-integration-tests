module bsg_ready_to_credit_flow_converter(clk_i, reset_i, v_i, ready_o, v_o, credit_i);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire [3:0] _16_;
  wire [3:0] _17_;
  input clk_i;
  wire clk_i;
  wire [3:0] credit_cnt;
  wire \credit_counter.clk_i ;
  reg [3:0] \credit_counter.count_o ;
  wire \credit_counter.down_i ;
  wire \credit_counter.reset_i ;
  wire \credit_counter.up_i ;
  input credit_i;
  wire credit_i;
  wire down;
  output ready_o;
  wire ready_o;
  input reset_i;
  wire reset_i;
  wire up;
  input v_i;
  wire v_i;
  output v_o;
  wire v_o;
  assign _00_ = ~(\credit_counter.count_o [0] | \credit_counter.count_o [1]);
  assign _01_ = \credit_counter.count_o [2] | \credit_counter.count_o [3];
  assign _02_ = _00_ & ~(_01_);
  assign ready_o = ~_02_;
  assign v_o = v_i & ~(_02_);
  assign _03_ = v_o & ~(credit_i);
  assign _04_ = _03_ ^ \credit_counter.count_o [1];
  assign _05_ = ~\credit_counter.count_o [0];
  assign _06_ = ~(v_o ^ credit_i);
  assign _07_ = _06_ | _05_;
  assign _17_[1] = ~(_07_ ^ _04_);
  assign _08_ = \credit_counter.count_o [2] ^ \credit_counter.count_o [1];
  assign _09_ = _03_ | \credit_counter.count_o [1];
  assign _10_ = _04_ & ~(_07_);
  assign _11_ = _09_ & ~(_10_);
  assign _17_[2] = _11_ ^ _08_;
  assign _12_ = \credit_counter.count_o [2] ^ \credit_counter.count_o [3];
  assign _13_ = \credit_counter.count_o [2] | ~(\credit_counter.count_o [1]);
  assign _14_ = ~(_11_ | _08_);
  assign _15_ = _13_ & ~(_14_);
  assign _17_[3] = _15_ ^ _12_;
  assign _16_[0] = _06_ ^ _05_;
  always @(posedge clk_i)
    if (reset_i) \credit_counter.count_o [0] <= 1'h0;
    else \credit_counter.count_o [0] <= _16_[0];
  always @(posedge clk_i)
    if (reset_i) \credit_counter.count_o [1] <= 1'h0;
    else \credit_counter.count_o [1] <= _17_[1];
  always @(posedge clk_i)
    if (reset_i) \credit_counter.count_o [2] <= 1'h0;
    else \credit_counter.count_o [2] <= _17_[2];
  always @(posedge clk_i)
    if (reset_i) \credit_counter.count_o [3] <= 1'h0;
    else \credit_counter.count_o [3] <= _17_[3];
  assign _17_[0] = _16_[0];
  assign credit_cnt = \credit_counter.count_o ;
  assign \credit_counter.clk_i  = clk_i;
  assign \credit_counter.down_i  = v_o;
  assign \credit_counter.reset_i  = reset_i;
  assign \credit_counter.up_i  = credit_i;
  assign down = v_o;
  assign up = credit_i;
endmodule
