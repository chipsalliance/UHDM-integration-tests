module bsg_reduce_segmented(i, o);
  input [15:0] i;
  wire [15:0] i;
  output o;
  wire o;
  assign o = 1'hx;
endmodule
