module bsg_scatter_gather(vec_i, fwd_o, fwd_datapath_o, bk_o, bk_datapath_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  output [7:0] bk_datapath_o;
  wire [7:0] bk_datapath_o;
  output [7:0] bk_o;
  wire [7:0] bk_o;
  output [7:0] fwd_datapath_o;
  wire [7:0] fwd_datapath_o;
  output [7:0] fwd_o;
  wire [7:0] fwd_o;
  input [3:0] vec_i;
  wire [3:0] vec_i;
  assign _00_ = ~vec_i[3];
  assign _01_ = ~vec_i[2];
  assign bk_o[2] = vec_i[0] | ~(vec_i[1]);
  assign _02_ = vec_i[2] ? bk_o[2] : vec_i[0];
  assign _03_ = _00_ & ~(_02_);
  assign _04_ = vec_i[3] & ~(_02_);
  assign fwd_o[0] = _04_ | _03_;
  assign fwd_o[1] = ~(vec_i[1] | vec_i[0]);
  assign _05_ = vec_i[1] | vec_i[0];
  assign bk_datapath_o[2] = vec_i[1] & vec_i[0];
  assign _06_ = bk_datapath_o[2] | ~(_05_);
  assign _07_ = _06_ | _01_;
  assign _08_ = vec_i[2] ? _06_ : _05_;
  assign fwd_o[2] = vec_i[3] ? _08_ : _07_;
  assign fwd_o[3] = ~(vec_i[1] & vec_i[0]);
  assign _09_ = fwd_o[3] | _01_;
  assign _10_ = vec_i[2] ? fwd_o[3] : bk_datapath_o[2];
  assign fwd_o[4] = vec_i[3] ? _10_ : _09_;
  assign _11_ = _05_ | _01_;
  assign fwd_o[5] = _11_ | _00_;
  assign _12_ = vec_i[1] & ~(vec_i[0]);
  assign _13_ = vec_i[2] & ~(_12_);
  assign fwd_o[6] = _13_ | _00_;
  assign _14_ = vec_i[2] & ~(bk_datapath_o[2]);
  assign fwd_o[7] = ~(_14_ & vec_i[3]);
  assign _15_ = ~(vec_i[1] ^ vec_i[0]);
  assign _16_ = _15_ | _01_;
  assign _17_ = _00_ & ~(_16_);
  assign _18_ = vec_i[3] & ~(_16_);
  assign bk_datapath_o[4] = _18_ | _17_;
  assign _19_ = _00_ & ~(_09_);
  assign _20_ = vec_i[3] & ~(_09_);
  assign bk_datapath_o[5] = _20_ | _19_;
  assign _21_ = vec_i[1] ^ vec_i[0];
  assign _22_ = vec_i[2] ? _06_ : _21_;
  assign bk_datapath_o[6] = _22_ & ~(_00_);
  assign _23_ = vec_i[2] ? _05_ : bk_datapath_o[2];
  assign bk_datapath_o[7] = _23_ & ~(_00_);
  assign _24_ = ~vec_i[0];
  assign _25_ = ~(_05_ & bk_o[2]);
  assign _26_ = vec_i[2] ? _24_ : _25_;
  assign bk_o[1] = vec_i[3] ? _24_ : _26_;
  assign _27_ = ~(vec_i[3] | vec_i[1]);
  assign _28_ = vec_i[3] & ~(vec_i[1]);
  assign bk_o[3] = _28_ | _27_;
  assign _29_ = _15_ & ~(_01_);
  assign _30_ = _00_ & ~(_29_);
  assign _31_ = vec_i[3] & ~(_29_);
  assign bk_o[4] = _31_ | _30_;
  assign _32_ = vec_i[3] & ~(_14_);
  assign _33_ = _00_ & ~(_14_);
  assign bk_o[5] = _33_ | _32_;
  assign bk_o[6] = _22_ | _00_;
  assign bk_o[7] = _23_ | _00_;
  assign _34_ = _12_ & ~(vec_i[3]);
  assign fwd_datapath_o[0] = _34_ | _04_;
  assign _35_ = vec_i[2] & ~(_05_);
  assign fwd_datapath_o[1] = vec_i[3] ? fwd_o[1] : _35_;
  assign _36_ = vec_i[2] ? _05_ : _15_;
  assign fwd_datapath_o[3] = vec_i[3] & ~(_36_);
  assign _37_ = vec_i[2] ? _15_ : fwd_o[3];
  assign fwd_datapath_o[4] = vec_i[3] & ~(_37_);
  assign { bk_datapath_o[3], bk_datapath_o[1:0] } = 3'h0;
  assign bk_o[0] = bk_o[1];
  assign { fwd_datapath_o[7:5], fwd_datapath_o[2] } = { 3'h0, bk_datapath_o[4] };
endmodule
