module top(output byte o);
   byte b[] = {1, 1, 1};
   assign o = b.and;
endmodule
