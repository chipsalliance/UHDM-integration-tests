module bsg_wait_cycles(clk_i, reset_i, activate_i, ready_r_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  input activate_i;
  wire activate_i;
  input clk_i;
  wire clk_i;
  wire [4:0] ctr_n;
  reg [4:0] ctr_r;
  output ready_r_o;
  reg ready_r_o;
  input reset_i;
  wire reset_i;
  assign _01_ = ctr_r[1] | ctr_r[0];
  assign _02_ = ctr_r[3] | ctr_r[2];
  assign _03_ = _02_ | _01_;
  assign _04_ = ctr_r[4] & ~(_03_);
  assign _05_ = ctr_r[3] & ctr_r[2];
  assign _06_ = ~(ctr_r[1] & ctr_r[0]);
  assign _07_ = _05_ & ~(_06_);
  assign _08_ = _07_ ^ ctr_r[4];
  assign _09_ = _04_ ? ctr_r[4] : _08_;
  assign _10_ = _09_ & ~(activate_i);
  assign ctr_n[4] = _10_ | reset_i;
  assign _11_ = ~reset_i;
  assign _12_ = _04_ ^ ctr_r[0];
  assign _13_ = _12_ | activate_i;
  assign ctr_n[0] = _11_ & ~(_13_);
  assign _14_ = ctr_r[1] ^ ctr_r[0];
  assign _15_ = _04_ ? ctr_r[1] : _14_;
  assign _16_ = activate_i | ~(_15_);
  assign ctr_n[1] = _11_ & ~(_16_);
  assign _17_ = ~ctr_r[2];
  assign _18_ = _06_ ^ ctr_r[2];
  assign _19_ = _04_ ? _17_ : _18_;
  assign _20_ = _19_ | activate_i;
  assign ctr_n[2] = _11_ & ~(_20_);
  assign _21_ = ctr_r[2] & ~(_06_);
  assign _22_ = _21_ ^ ctr_r[3];
  assign _23_ = _04_ ? ctr_r[3] : _22_;
  assign _24_ = activate_i | ~(_23_);
  assign ctr_n[3] = _11_ & ~(_24_);
  assign _25_ = ctr_n[1] | ctr_n[0];
  assign _26_ = ctr_n[3] | ctr_n[2];
  assign _27_ = _26_ | _25_;
  assign _00_ = ctr_n[4] & ~(_27_);
  always @(posedge clk_i)
    ready_r_o <= _00_;
  always @(posedge clk_i)
    ctr_r[0] <= ctr_n[0];
  always @(posedge clk_i)
    ctr_r[1] <= ctr_n[1];
  always @(posedge clk_i)
    ctr_r[2] <= ctr_n[2];
  always @(posedge clk_i)
    ctr_r[3] <= ctr_n[3];
  always @(posedge clk_i)
    ctr_r[4] <= ctr_n[4];
endmodule
