module bsg_flow_counter(clk_i, reset_i, v_i, ready_i, yumi_i, count_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire [6:0] _31_;
  wire [6:0] _32_;
  input clk_i;
  wire clk_i;
  output [6:0] count_o;
  wire [6:0] count_o;
  wire enque;
  wire \gen_blk_0.counter.clk_i ;
  reg [6:0] \gen_blk_0.counter.count_o ;
  wire \gen_blk_0.counter.down_i ;
  wire \gen_blk_0.counter.reset_i ;
  wire \gen_blk_0.counter.up_i ;
  input ready_i;
  wire ready_i;
  input reset_i;
  wire reset_i;
  input v_i;
  wire v_i;
  input yumi_i;
  wire yumi_i;
  assign _00_ = yumi_i & ~(\gen_blk_0.counter.count_o [0]);
  assign _01_ = _00_ ^ \gen_blk_0.counter.count_o [1];
  assign _02_ = ~(yumi_i ^ \gen_blk_0.counter.count_o [0]);
  assign _03_ = ~(ready_i & v_i);
  assign _04_ = _03_ | _02_;
  assign _32_[1] = ~(_04_ ^ _01_);
  assign _05_ = \gen_blk_0.counter.count_o [2] ^ \gen_blk_0.counter.count_o [1];
  assign _06_ = _00_ | \gen_blk_0.counter.count_o [1];
  assign _07_ = _01_ & ~(_04_);
  assign _08_ = _07_ | ~(_06_);
  assign _32_[2] = ~(_08_ ^ _05_);
  assign _09_ = \gen_blk_0.counter.count_o [2] ^ \gen_blk_0.counter.count_o [3];
  assign _10_ = \gen_blk_0.counter.count_o [2] | ~(\gen_blk_0.counter.count_o [1]);
  assign _11_ = _08_ & ~(_05_);
  assign _12_ = _10_ & ~(_11_);
  assign _32_[3] = _12_ ^ _09_;
  assign _13_ = \gen_blk_0.counter.count_o [3] ^ \gen_blk_0.counter.count_o [4];
  assign _14_ = \gen_blk_0.counter.count_o [3] | ~(\gen_blk_0.counter.count_o [2]);
  assign _15_ = ~(_10_ | _09_);
  assign _16_ = _14_ & ~(_15_);
  assign _17_ = _09_ | _05_;
  assign _18_ = _08_ & ~(_17_);
  assign _19_ = _16_ & ~(_18_);
  assign _32_[4] = _19_ ^ _13_;
  assign _20_ = \gen_blk_0.counter.count_o [4] ^ \gen_blk_0.counter.count_o [5];
  assign _21_ = \gen_blk_0.counter.count_o [4] | ~(\gen_blk_0.counter.count_o [3]);
  assign _22_ = ~(_19_ | _13_);
  assign _23_ = _21_ & ~(_22_);
  assign _32_[5] = _23_ ^ _20_;
  assign _24_ = \gen_blk_0.counter.count_o [5] ^ \gen_blk_0.counter.count_o [6];
  assign _25_ = \gen_blk_0.counter.count_o [5] | ~(\gen_blk_0.counter.count_o [4]);
  assign _26_ = ~(_21_ | _20_);
  assign _27_ = _25_ & ~(_26_);
  assign _28_ = _20_ | _13_;
  assign _29_ = ~(_28_ | _19_);
  assign _30_ = _27_ & ~(_29_);
  assign _32_[6] = _30_ ^ _24_;
  assign _31_[0] = _03_ ^ _02_;
  always @(posedge clk_i)
    if (reset_i) \gen_blk_0.counter.count_o [0] <= 1'h0;
    else \gen_blk_0.counter.count_o [0] <= _31_[0];
  always @(posedge clk_i)
    if (reset_i) \gen_blk_0.counter.count_o [1] <= 1'h0;
    else \gen_blk_0.counter.count_o [1] <= _32_[1];
  always @(posedge clk_i)
    if (reset_i) \gen_blk_0.counter.count_o [2] <= 1'h0;
    else \gen_blk_0.counter.count_o [2] <= _32_[2];
  always @(posedge clk_i)
    if (reset_i) \gen_blk_0.counter.count_o [3] <= 1'h0;
    else \gen_blk_0.counter.count_o [3] <= _32_[3];
  always @(posedge clk_i)
    if (reset_i) \gen_blk_0.counter.count_o [4] <= 1'h0;
    else \gen_blk_0.counter.count_o [4] <= _32_[4];
  always @(posedge clk_i)
    if (reset_i) \gen_blk_0.counter.count_o [5] <= 1'h0;
    else \gen_blk_0.counter.count_o [5] <= _32_[5];
  always @(posedge clk_i)
    if (reset_i) \gen_blk_0.counter.count_o [6] <= 1'h0;
    else \gen_blk_0.counter.count_o [6] <= _32_[6];
  assign _32_[0] = _31_[0];
  assign count_o = \gen_blk_0.counter.count_o ;
  assign enque = \gen_blk_0.counter.up_i ;
  assign \gen_blk_0.counter.clk_i  = clk_i;
  assign \gen_blk_0.counter.down_i  = yumi_i;
  assign \gen_blk_0.counter.reset_i  = reset_i;
endmodule
