module bsg_cache_decode(opcode_i, decode_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  output [20:0] decode_o;
  wire [20:0] decode_o;
  input [5:0] opcode_i;
  wire [5:0] opcode_i;
  assign _008_ = opcode_i[1] | opcode_i[0];
  assign _009_ = opcode_i[3] | opcode_i[2];
  assign _010_ = ~(_009_ | _008_);
  assign _011_ = opcode_i[4] & ~(opcode_i[5]);
  assign decode_o[14] = _011_ & _010_;
  assign decode_o[5] = ~decode_o[14];
  assign _012_ = opcode_i[1] | ~(opcode_i[0]);
  assign _013_ = ~(_012_ | _009_);
  assign decode_o[13] = _013_ & _011_;
  assign _014_ = opcode_i[0] | ~(opcode_i[1]);
  assign _015_ = ~(_014_ | _009_);
  assign decode_o[12] = _015_ & _011_;
  assign _016_ = ~(opcode_i[1] & opcode_i[0]);
  assign _017_ = ~(_016_ | _009_);
  assign decode_o[11] = _017_ & _011_;
  assign _018_ = opcode_i[2] | ~(opcode_i[3]);
  assign _019_ = ~(_018_ | _008_);
  assign decode_o[10] = _019_ & _011_;
  assign _020_ = ~(_018_ | _012_);
  assign decode_o[9] = _020_ & _011_;
  assign _021_ = ~(_018_ | _014_);
  assign decode_o[8] = _021_ & _011_;
  assign _022_ = ~(_018_ | _016_);
  assign decode_o[7] = _022_ & _011_;
  assign _023_ = ~(opcode_i[3] & opcode_i[2]);
  assign _024_ = ~(_023_ | _008_);
  assign decode_o[6] = _024_ & _011_;
  assign _025_ = ~(_008_ | opcode_i[2]);
  assign _026_ = opcode_i[3] & ~(_025_);
  assign decode_o[4] = opcode_i[5] & ~(_026_);
  assign _027_ = opcode_i[5] | opcode_i[4];
  assign _028_ = _010_ & ~(_027_);
  assign _029_ = _013_ & ~(_027_);
  assign _030_ = _029_ | _028_;
  assign _031_ = _015_ & ~(_027_);
  assign _032_ = _031_ | _030_;
  assign _033_ = _017_ & ~(_027_);
  assign _034_ = _033_ | _032_;
  assign decode_o[18] = _034_ | decode_o[4];
  assign _035_ = opcode_i[3] | ~(opcode_i[2]);
  assign _036_ = _035_ | _008_;
  assign _037_ = ~(_036_ | _027_);
  assign _038_ = _037_ | _034_;
  assign _039_ = _035_ | _012_;
  assign _040_ = ~(_039_ | _027_);
  assign _041_ = _040_ | _038_;
  assign _042_ = _035_ | _014_;
  assign _043_ = ~(_042_ | _027_);
  assign _044_ = _043_ | _041_;
  assign _045_ = _035_ | _016_;
  assign _046_ = ~(_045_ | _027_);
  assign _047_ = _046_ | _044_;
  assign _048_ = _024_ & ~(_027_);
  assign decode_o[16] = _048_ | _047_;
  assign _049_ = _019_ & ~(_027_);
  assign _050_ = _020_ & ~(_027_);
  assign _051_ = _050_ | _049_;
  assign _052_ = _021_ & ~(_027_);
  assign _053_ = _052_ | _051_;
  assign _054_ = _022_ & ~(_027_);
  assign _055_ = _054_ | _053_;
  assign _056_ = _023_ | _012_;
  assign _057_ = ~(_056_ | _027_);
  assign decode_o[15] = _057_ | _055_;
  assign _058_ = opcode_i[3] | ~(opcode_i[0]);
  assign decode_o[0] = opcode_i[5] & ~(_058_);
  assign _059_ = opcode_i[3] | ~(opcode_i[1]);
  assign decode_o[1] = opcode_i[5] & ~(_059_);
  assign decode_o[2] = opcode_i[5] & ~(_035_);
  assign _060_ = ~(_025_ & opcode_i[3]);
  assign decode_o[3] = opcode_i[5] & ~(_060_);
  assign _000_ = opcode_i[0] & ~(opcode_i[2]);
  assign _001_ = opcode_i[3] ? _000_ : opcode_i[0];
  assign _002_ = _001_ & ~(opcode_i[4]);
  assign _003_ = opcode_i[4] & ~(_026_);
  assign decode_o[19] = opcode_i[5] ? _003_ : _002_;
  assign _004_ = ~_026_;
  assign _005_ = opcode_i[1] & ~(opcode_i[2]);
  assign _006_ = opcode_i[3] ? _005_ : opcode_i[1];
  assign _007_ = _006_ & ~(opcode_i[4]);
  assign decode_o[20] = opcode_i[5] ? _004_ : _007_;
  assign decode_o[17] = _057_ | _048_;
endmodule
