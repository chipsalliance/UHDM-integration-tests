module bsg_fifo_shift_datapath(clk_i, data_i, sel_i, data_o);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  input clk_i;
  wire clk_i;
  input [15:0] data_i;
  wire [15:0] data_i;
  output [15:0] data_o;
  reg [15:0] data_o;
  wire [511:0] r;
  wire [511:0] r_n;
  input [63:0] sel_i;
  wire [63:0] sel_i;
  assign _0007_ = sel_i[14] ^ sel_i[15];
  assign _0006_ = sel_i[12] ^ sel_i[13];
  assign _0005_ = sel_i[10] ^ sel_i[11];
  assign _0004_ = sel_i[8] ^ sel_i[9];
  assign _0003_ = sel_i[6] ^ sel_i[7];
  assign _0002_ = sel_i[4] ^ sel_i[5];
  assign _0001_ = sel_i[2] ^ sel_i[3];
  assign _0000_ = sel_i[0] ^ sel_i[1];
  assign _0031_ = sel_i[62] ^ sel_i[63];
  assign _0030_ = sel_i[60] ^ sel_i[61];
  assign _0029_ = sel_i[58] ^ sel_i[59];
  assign _0028_ = sel_i[56] ^ sel_i[57];
  assign _0027_ = sel_i[54] ^ sel_i[55];
  assign _0026_ = sel_i[52] ^ sel_i[53];
  assign _0025_ = sel_i[50] ^ sel_i[51];
  assign _0024_ = sel_i[48] ^ sel_i[49];
  assign _0023_ = sel_i[46] ^ sel_i[47];
  assign _0022_ = sel_i[44] ^ sel_i[45];
  assign _0021_ = sel_i[42] ^ sel_i[43];
  assign _0020_ = sel_i[40] ^ sel_i[41];
  assign _0019_ = sel_i[38] ^ sel_i[39];
  assign _0018_ = sel_i[36] ^ sel_i[37];
  assign _0017_ = sel_i[34] ^ sel_i[35];
  assign _0016_ = sel_i[32] ^ sel_i[33];
  assign _0015_ = sel_i[30] ^ sel_i[31];
  assign _0032_ = sel_i[62] | ~(sel_i[63]);
  assign _0014_ = sel_i[28] ^ sel_i[29];
  assign _0013_ = sel_i[26] ^ sel_i[27];
  assign _0012_ = sel_i[24] ^ sel_i[25];
  assign _0011_ = sel_i[22] ^ sel_i[23];
  assign _0010_ = sel_i[20] ^ sel_i[21];
  assign _0009_ = sel_i[18] ^ sel_i[19];
  assign _0008_ = sel_i[16] ^ sel_i[17];
  assign _0033_ = sel_i[33] & ~(sel_i[32]);
  assign r_n[256] = _0033_ ? data_i[0] : r[272];
  assign r_n[257] = _0033_ ? data_i[1] : r[273];
  assign r_n[258] = _0033_ ? data_i[2] : r[274];
  assign r_n[259] = _0033_ ? data_i[3] : r[275];
  assign r_n[260] = _0033_ ? data_i[4] : r[276];
  assign r_n[261] = _0033_ ? data_i[5] : r[277];
  assign r_n[262] = _0033_ ? data_i[6] : r[278];
  assign r_n[263] = _0033_ ? data_i[7] : r[279];
  assign r_n[264] = _0033_ ? data_i[8] : r[280];
  assign r_n[265] = _0033_ ? data_i[9] : r[281];
  assign r_n[266] = _0033_ ? data_i[10] : r[282];
  assign r_n[267] = _0033_ ? data_i[11] : r[283];
  assign r_n[268] = _0033_ ? data_i[12] : r[284];
  assign r_n[269] = _0033_ ? data_i[13] : r[285];
  assign r_n[270] = _0033_ ? data_i[14] : r[286];
  assign r_n[271] = _0033_ ? data_i[15] : r[287];
  assign _0034_ = sel_i[31] & ~(sel_i[30]);
  assign r_n[240] = _0034_ ? data_i[0] : r[256];
  assign r_n[241] = _0034_ ? data_i[1] : r[257];
  assign r_n[242] = _0034_ ? data_i[2] : r[258];
  assign r_n[243] = _0034_ ? data_i[3] : r[259];
  assign r_n[244] = _0034_ ? data_i[4] : r[260];
  assign r_n[245] = _0034_ ? data_i[5] : r[261];
  assign r_n[246] = _0034_ ? data_i[6] : r[262];
  assign r_n[247] = _0034_ ? data_i[7] : r[263];
  assign r_n[248] = _0034_ ? data_i[8] : r[264];
  assign r_n[249] = _0034_ ? data_i[9] : r[265];
  assign r_n[250] = _0034_ ? data_i[10] : r[266];
  assign r_n[251] = _0034_ ? data_i[11] : r[267];
  assign r_n[252] = _0034_ ? data_i[12] : r[268];
  assign r_n[253] = _0034_ ? data_i[13] : r[269];
  assign r_n[254] = _0034_ ? data_i[14] : r[270];
  assign r_n[255] = _0034_ ? data_i[15] : r[271];
  assign _0035_ = sel_i[29] & ~(sel_i[28]);
  assign r_n[224] = _0035_ ? data_i[0] : r[240];
  assign r_n[225] = _0035_ ? data_i[1] : r[241];
  assign r_n[226] = _0035_ ? data_i[2] : r[242];
  assign r_n[227] = _0035_ ? data_i[3] : r[243];
  assign r_n[228] = _0035_ ? data_i[4] : r[244];
  assign r_n[229] = _0035_ ? data_i[5] : r[245];
  assign r_n[230] = _0035_ ? data_i[6] : r[246];
  assign r_n[231] = _0035_ ? data_i[7] : r[247];
  assign r_n[232] = _0035_ ? data_i[8] : r[248];
  assign r_n[233] = _0035_ ? data_i[9] : r[249];
  assign r_n[234] = _0035_ ? data_i[10] : r[250];
  assign r_n[235] = _0035_ ? data_i[11] : r[251];
  assign r_n[236] = _0035_ ? data_i[12] : r[252];
  assign r_n[237] = _0035_ ? data_i[13] : r[253];
  assign r_n[238] = _0035_ ? data_i[14] : r[254];
  assign r_n[239] = _0035_ ? data_i[15] : r[255];
  assign _0036_ = sel_i[27] & ~(sel_i[26]);
  assign r_n[208] = _0036_ ? data_i[0] : r[224];
  assign r_n[209] = _0036_ ? data_i[1] : r[225];
  assign r_n[210] = _0036_ ? data_i[2] : r[226];
  assign r_n[211] = _0036_ ? data_i[3] : r[227];
  assign r_n[212] = _0036_ ? data_i[4] : r[228];
  assign r_n[213] = _0036_ ? data_i[5] : r[229];
  assign r_n[214] = _0036_ ? data_i[6] : r[230];
  assign r_n[215] = _0036_ ? data_i[7] : r[231];
  assign r_n[216] = _0036_ ? data_i[8] : r[232];
  assign r_n[217] = _0036_ ? data_i[9] : r[233];
  assign r_n[218] = _0036_ ? data_i[10] : r[234];
  assign r_n[219] = _0036_ ? data_i[11] : r[235];
  assign r_n[220] = _0036_ ? data_i[12] : r[236];
  assign r_n[221] = _0036_ ? data_i[13] : r[237];
  assign r_n[222] = _0036_ ? data_i[14] : r[238];
  assign r_n[223] = _0036_ ? data_i[15] : r[239];
  assign _0037_ = sel_i[25] & ~(sel_i[24]);
  assign r_n[192] = _0037_ ? data_i[0] : r[208];
  assign r_n[193] = _0037_ ? data_i[1] : r[209];
  assign r_n[194] = _0037_ ? data_i[2] : r[210];
  assign r_n[195] = _0037_ ? data_i[3] : r[211];
  assign r_n[196] = _0037_ ? data_i[4] : r[212];
  assign r_n[197] = _0037_ ? data_i[5] : r[213];
  assign r_n[198] = _0037_ ? data_i[6] : r[214];
  assign r_n[199] = _0037_ ? data_i[7] : r[215];
  assign r_n[200] = _0037_ ? data_i[8] : r[216];
  assign r_n[201] = _0037_ ? data_i[9] : r[217];
  assign r_n[202] = _0037_ ? data_i[10] : r[218];
  assign r_n[203] = _0037_ ? data_i[11] : r[219];
  assign r_n[204] = _0037_ ? data_i[12] : r[220];
  assign r_n[205] = _0037_ ? data_i[13] : r[221];
  assign r_n[206] = _0037_ ? data_i[14] : r[222];
  assign r_n[207] = _0037_ ? data_i[15] : r[223];
  assign _0038_ = sel_i[23] & ~(sel_i[22]);
  assign r_n[176] = _0038_ ? data_i[0] : r[192];
  assign r_n[177] = _0038_ ? data_i[1] : r[193];
  assign r_n[178] = _0038_ ? data_i[2] : r[194];
  assign r_n[179] = _0038_ ? data_i[3] : r[195];
  assign r_n[180] = _0038_ ? data_i[4] : r[196];
  assign r_n[181] = _0038_ ? data_i[5] : r[197];
  assign r_n[182] = _0038_ ? data_i[6] : r[198];
  assign r_n[183] = _0038_ ? data_i[7] : r[199];
  assign r_n[184] = _0038_ ? data_i[8] : r[200];
  assign r_n[185] = _0038_ ? data_i[9] : r[201];
  assign r_n[186] = _0038_ ? data_i[10] : r[202];
  assign r_n[187] = _0038_ ? data_i[11] : r[203];
  assign r_n[188] = _0038_ ? data_i[12] : r[204];
  assign r_n[189] = _0038_ ? data_i[13] : r[205];
  assign r_n[190] = _0038_ ? data_i[14] : r[206];
  assign r_n[191] = _0038_ ? data_i[15] : r[207];
  assign _0039_ = sel_i[21] & ~(sel_i[20]);
  assign r_n[160] = _0039_ ? data_i[0] : r[176];
  assign r_n[161] = _0039_ ? data_i[1] : r[177];
  assign r_n[162] = _0039_ ? data_i[2] : r[178];
  assign r_n[163] = _0039_ ? data_i[3] : r[179];
  assign r_n[164] = _0039_ ? data_i[4] : r[180];
  assign r_n[165] = _0039_ ? data_i[5] : r[181];
  assign r_n[166] = _0039_ ? data_i[6] : r[182];
  assign r_n[167] = _0039_ ? data_i[7] : r[183];
  assign r_n[168] = _0039_ ? data_i[8] : r[184];
  assign r_n[169] = _0039_ ? data_i[9] : r[185];
  assign r_n[170] = _0039_ ? data_i[10] : r[186];
  assign r_n[171] = _0039_ ? data_i[11] : r[187];
  assign r_n[172] = _0039_ ? data_i[12] : r[188];
  assign r_n[173] = _0039_ ? data_i[13] : r[189];
  assign r_n[174] = _0039_ ? data_i[14] : r[190];
  assign r_n[175] = _0039_ ? data_i[15] : r[191];
  assign _0040_ = sel_i[19] & ~(sel_i[18]);
  assign r_n[144] = _0040_ ? data_i[0] : r[160];
  assign r_n[145] = _0040_ ? data_i[1] : r[161];
  assign r_n[146] = _0040_ ? data_i[2] : r[162];
  assign r_n[147] = _0040_ ? data_i[3] : r[163];
  assign r_n[148] = _0040_ ? data_i[4] : r[164];
  assign r_n[149] = _0040_ ? data_i[5] : r[165];
  assign r_n[150] = _0040_ ? data_i[6] : r[166];
  assign r_n[151] = _0040_ ? data_i[7] : r[167];
  assign r_n[152] = _0040_ ? data_i[8] : r[168];
  assign r_n[153] = _0040_ ? data_i[9] : r[169];
  assign r_n[154] = _0040_ ? data_i[10] : r[170];
  assign r_n[155] = _0040_ ? data_i[11] : r[171];
  assign r_n[156] = _0040_ ? data_i[12] : r[172];
  assign r_n[157] = _0040_ ? data_i[13] : r[173];
  assign r_n[158] = _0040_ ? data_i[14] : r[174];
  assign r_n[159] = _0040_ ? data_i[15] : r[175];
  assign _0041_ = sel_i[17] & ~(sel_i[16]);
  assign r_n[128] = _0041_ ? data_i[0] : r[144];
  assign r_n[129] = _0041_ ? data_i[1] : r[145];
  assign r_n[130] = _0041_ ? data_i[2] : r[146];
  assign r_n[131] = _0041_ ? data_i[3] : r[147];
  assign r_n[132] = _0041_ ? data_i[4] : r[148];
  assign r_n[133] = _0041_ ? data_i[5] : r[149];
  assign r_n[134] = _0041_ ? data_i[6] : r[150];
  assign r_n[135] = _0041_ ? data_i[7] : r[151];
  assign r_n[136] = _0041_ ? data_i[8] : r[152];
  assign r_n[137] = _0041_ ? data_i[9] : r[153];
  assign r_n[138] = _0041_ ? data_i[10] : r[154];
  assign r_n[139] = _0041_ ? data_i[11] : r[155];
  assign r_n[140] = _0041_ ? data_i[12] : r[156];
  assign r_n[141] = _0041_ ? data_i[13] : r[157];
  assign r_n[142] = _0041_ ? data_i[14] : r[158];
  assign r_n[143] = _0041_ ? data_i[15] : r[159];
  assign _0042_ = sel_i[15] & ~(sel_i[14]);
  assign r_n[112] = _0042_ ? data_i[0] : r[128];
  assign r_n[113] = _0042_ ? data_i[1] : r[129];
  assign r_n[114] = _0042_ ? data_i[2] : r[130];
  assign r_n[115] = _0042_ ? data_i[3] : r[131];
  assign r_n[116] = _0042_ ? data_i[4] : r[132];
  assign r_n[117] = _0042_ ? data_i[5] : r[133];
  assign r_n[118] = _0042_ ? data_i[6] : r[134];
  assign r_n[119] = _0042_ ? data_i[7] : r[135];
  assign r_n[120] = _0042_ ? data_i[8] : r[136];
  assign r_n[121] = _0042_ ? data_i[9] : r[137];
  assign r_n[122] = _0042_ ? data_i[10] : r[138];
  assign r_n[123] = _0042_ ? data_i[11] : r[139];
  assign r_n[124] = _0042_ ? data_i[12] : r[140];
  assign r_n[125] = _0042_ ? data_i[13] : r[141];
  assign r_n[126] = _0042_ ? data_i[14] : r[142];
  assign r_n[127] = _0042_ ? data_i[15] : r[143];
  assign _0043_ = sel_i[13] & ~(sel_i[12]);
  assign r_n[96] = _0043_ ? data_i[0] : r[112];
  assign r_n[97] = _0043_ ? data_i[1] : r[113];
  assign r_n[98] = _0043_ ? data_i[2] : r[114];
  assign r_n[99] = _0043_ ? data_i[3] : r[115];
  assign r_n[100] = _0043_ ? data_i[4] : r[116];
  assign r_n[101] = _0043_ ? data_i[5] : r[117];
  assign r_n[102] = _0043_ ? data_i[6] : r[118];
  assign r_n[103] = _0043_ ? data_i[7] : r[119];
  assign r_n[104] = _0043_ ? data_i[8] : r[120];
  assign r_n[105] = _0043_ ? data_i[9] : r[121];
  assign r_n[106] = _0043_ ? data_i[10] : r[122];
  assign r_n[107] = _0043_ ? data_i[11] : r[123];
  assign r_n[108] = _0043_ ? data_i[12] : r[124];
  assign r_n[109] = _0043_ ? data_i[13] : r[125];
  assign r_n[110] = _0043_ ? data_i[14] : r[126];
  assign r_n[111] = _0043_ ? data_i[15] : r[127];
  assign _0044_ = sel_i[11] & ~(sel_i[10]);
  assign r_n[80] = _0044_ ? data_i[0] : r[96];
  assign r_n[81] = _0044_ ? data_i[1] : r[97];
  assign r_n[82] = _0044_ ? data_i[2] : r[98];
  assign r_n[83] = _0044_ ? data_i[3] : r[99];
  assign r_n[84] = _0044_ ? data_i[4] : r[100];
  assign r_n[85] = _0044_ ? data_i[5] : r[101];
  assign r_n[86] = _0044_ ? data_i[6] : r[102];
  assign r_n[87] = _0044_ ? data_i[7] : r[103];
  assign r_n[88] = _0044_ ? data_i[8] : r[104];
  assign r_n[89] = _0044_ ? data_i[9] : r[105];
  assign r_n[90] = _0044_ ? data_i[10] : r[106];
  assign r_n[91] = _0044_ ? data_i[11] : r[107];
  assign r_n[92] = _0044_ ? data_i[12] : r[108];
  assign r_n[93] = _0044_ ? data_i[13] : r[109];
  assign r_n[94] = _0044_ ? data_i[14] : r[110];
  assign r_n[95] = _0044_ ? data_i[15] : r[111];
  assign _0045_ = sel_i[9] & ~(sel_i[8]);
  assign r_n[64] = _0045_ ? data_i[0] : r[80];
  assign r_n[65] = _0045_ ? data_i[1] : r[81];
  assign r_n[66] = _0045_ ? data_i[2] : r[82];
  assign r_n[67] = _0045_ ? data_i[3] : r[83];
  assign r_n[68] = _0045_ ? data_i[4] : r[84];
  assign r_n[69] = _0045_ ? data_i[5] : r[85];
  assign r_n[70] = _0045_ ? data_i[6] : r[86];
  assign r_n[71] = _0045_ ? data_i[7] : r[87];
  assign r_n[72] = _0045_ ? data_i[8] : r[88];
  assign r_n[73] = _0045_ ? data_i[9] : r[89];
  assign r_n[74] = _0045_ ? data_i[10] : r[90];
  assign r_n[75] = _0045_ ? data_i[11] : r[91];
  assign r_n[76] = _0045_ ? data_i[12] : r[92];
  assign r_n[77] = _0045_ ? data_i[13] : r[93];
  assign r_n[78] = _0045_ ? data_i[14] : r[94];
  assign r_n[79] = _0045_ ? data_i[15] : r[95];
  assign _0046_ = sel_i[7] & ~(sel_i[6]);
  assign r_n[48] = _0046_ ? data_i[0] : r[64];
  assign r_n[49] = _0046_ ? data_i[1] : r[65];
  assign r_n[50] = _0046_ ? data_i[2] : r[66];
  assign r_n[51] = _0046_ ? data_i[3] : r[67];
  assign r_n[52] = _0046_ ? data_i[4] : r[68];
  assign r_n[53] = _0046_ ? data_i[5] : r[69];
  assign r_n[54] = _0046_ ? data_i[6] : r[70];
  assign r_n[55] = _0046_ ? data_i[7] : r[71];
  assign r_n[56] = _0046_ ? data_i[8] : r[72];
  assign r_n[57] = _0046_ ? data_i[9] : r[73];
  assign r_n[58] = _0046_ ? data_i[10] : r[74];
  assign r_n[59] = _0046_ ? data_i[11] : r[75];
  assign r_n[60] = _0046_ ? data_i[12] : r[76];
  assign r_n[61] = _0046_ ? data_i[13] : r[77];
  assign r_n[62] = _0046_ ? data_i[14] : r[78];
  assign r_n[63] = _0046_ ? data_i[15] : r[79];
  assign _0047_ = sel_i[5] & ~(sel_i[4]);
  assign r_n[32] = _0047_ ? data_i[0] : r[48];
  assign r_n[33] = _0047_ ? data_i[1] : r[49];
  assign r_n[34] = _0047_ ? data_i[2] : r[50];
  assign r_n[35] = _0047_ ? data_i[3] : r[51];
  assign r_n[36] = _0047_ ? data_i[4] : r[52];
  assign r_n[37] = _0047_ ? data_i[5] : r[53];
  assign r_n[38] = _0047_ ? data_i[6] : r[54];
  assign r_n[39] = _0047_ ? data_i[7] : r[55];
  assign r_n[40] = _0047_ ? data_i[8] : r[56];
  assign r_n[41] = _0047_ ? data_i[9] : r[57];
  assign r_n[42] = _0047_ ? data_i[10] : r[58];
  assign r_n[43] = _0047_ ? data_i[11] : r[59];
  assign r_n[44] = _0047_ ? data_i[12] : r[60];
  assign r_n[45] = _0047_ ? data_i[13] : r[61];
  assign r_n[46] = _0047_ ? data_i[14] : r[62];
  assign r_n[47] = _0047_ ? data_i[15] : r[63];
  assign _0048_ = sel_i[3] & ~(sel_i[2]);
  assign r_n[16] = _0048_ ? data_i[0] : r[32];
  assign r_n[17] = _0048_ ? data_i[1] : r[33];
  assign r_n[18] = _0048_ ? data_i[2] : r[34];
  assign r_n[19] = _0048_ ? data_i[3] : r[35];
  assign r_n[20] = _0048_ ? data_i[4] : r[36];
  assign r_n[21] = _0048_ ? data_i[5] : r[37];
  assign r_n[22] = _0048_ ? data_i[6] : r[38];
  assign r_n[23] = _0048_ ? data_i[7] : r[39];
  assign r_n[24] = _0048_ ? data_i[8] : r[40];
  assign r_n[25] = _0048_ ? data_i[9] : r[41];
  assign r_n[26] = _0048_ ? data_i[10] : r[42];
  assign r_n[27] = _0048_ ? data_i[11] : r[43];
  assign r_n[28] = _0048_ ? data_i[12] : r[44];
  assign r_n[29] = _0048_ ? data_i[13] : r[45];
  assign r_n[30] = _0048_ ? data_i[14] : r[46];
  assign r_n[31] = _0048_ ? data_i[15] : r[47];
  assign _0049_ = sel_i[1] & ~(sel_i[0]);
  assign r_n[0] = _0049_ ? data_i[0] : r[16];
  assign r_n[1] = _0049_ ? data_i[1] : r[17];
  assign r_n[2] = _0049_ ? data_i[2] : r[18];
  assign r_n[3] = _0049_ ? data_i[3] : r[19];
  assign r_n[4] = _0049_ ? data_i[4] : r[20];
  assign r_n[5] = _0049_ ? data_i[5] : r[21];
  assign r_n[6] = _0049_ ? data_i[6] : r[22];
  assign r_n[7] = _0049_ ? data_i[7] : r[23];
  assign r_n[8] = _0049_ ? data_i[8] : r[24];
  assign r_n[9] = _0049_ ? data_i[9] : r[25];
  assign r_n[10] = _0049_ ? data_i[10] : r[26];
  assign r_n[11] = _0049_ ? data_i[11] : r[27];
  assign r_n[12] = _0049_ ? data_i[12] : r[28];
  assign r_n[13] = _0049_ ? data_i[13] : r[29];
  assign r_n[14] = _0049_ ? data_i[14] : r[30];
  assign r_n[15] = _0049_ ? data_i[15] : r[31];
  assign _0050_ = sel_i[61] & ~(sel_i[60]);
  assign r_n[480] = _0050_ ? data_i[0] : r[496];
  assign r_n[481] = _0050_ ? data_i[1] : r[497];
  assign r_n[482] = _0050_ ? data_i[2] : r[498];
  assign r_n[483] = _0050_ ? data_i[3] : r[499];
  assign r_n[484] = _0050_ ? data_i[4] : r[500];
  assign r_n[485] = _0050_ ? data_i[5] : r[501];
  assign r_n[486] = _0050_ ? data_i[6] : r[502];
  assign r_n[487] = _0050_ ? data_i[7] : r[503];
  assign r_n[488] = _0050_ ? data_i[8] : r[504];
  assign r_n[489] = _0050_ ? data_i[9] : r[505];
  assign r_n[490] = _0050_ ? data_i[10] : r[506];
  assign r_n[491] = _0050_ ? data_i[11] : r[507];
  assign r_n[492] = _0050_ ? data_i[12] : r[508];
  assign r_n[493] = _0050_ ? data_i[13] : r[509];
  assign r_n[494] = _0050_ ? data_i[14] : r[510];
  assign r_n[495] = _0050_ ? data_i[15] : r[511];
  assign _0051_ = sel_i[59] & ~(sel_i[58]);
  assign r_n[464] = _0051_ ? data_i[0] : r[480];
  assign r_n[465] = _0051_ ? data_i[1] : r[481];
  assign r_n[466] = _0051_ ? data_i[2] : r[482];
  assign r_n[467] = _0051_ ? data_i[3] : r[483];
  assign r_n[468] = _0051_ ? data_i[4] : r[484];
  assign r_n[469] = _0051_ ? data_i[5] : r[485];
  assign r_n[470] = _0051_ ? data_i[6] : r[486];
  assign r_n[471] = _0051_ ? data_i[7] : r[487];
  assign r_n[472] = _0051_ ? data_i[8] : r[488];
  assign r_n[473] = _0051_ ? data_i[9] : r[489];
  assign r_n[474] = _0051_ ? data_i[10] : r[490];
  assign r_n[475] = _0051_ ? data_i[11] : r[491];
  assign r_n[476] = _0051_ ? data_i[12] : r[492];
  assign r_n[477] = _0051_ ? data_i[13] : r[493];
  assign r_n[478] = _0051_ ? data_i[14] : r[494];
  assign r_n[479] = _0051_ ? data_i[15] : r[495];
  assign _0052_ = sel_i[57] & ~(sel_i[56]);
  assign r_n[448] = _0052_ ? data_i[0] : r[464];
  assign r_n[449] = _0052_ ? data_i[1] : r[465];
  assign r_n[450] = _0052_ ? data_i[2] : r[466];
  assign r_n[451] = _0052_ ? data_i[3] : r[467];
  assign r_n[452] = _0052_ ? data_i[4] : r[468];
  assign r_n[453] = _0052_ ? data_i[5] : r[469];
  assign r_n[454] = _0052_ ? data_i[6] : r[470];
  assign r_n[455] = _0052_ ? data_i[7] : r[471];
  assign r_n[456] = _0052_ ? data_i[8] : r[472];
  assign r_n[457] = _0052_ ? data_i[9] : r[473];
  assign r_n[458] = _0052_ ? data_i[10] : r[474];
  assign r_n[459] = _0052_ ? data_i[11] : r[475];
  assign r_n[460] = _0052_ ? data_i[12] : r[476];
  assign r_n[461] = _0052_ ? data_i[13] : r[477];
  assign r_n[462] = _0052_ ? data_i[14] : r[478];
  assign r_n[463] = _0052_ ? data_i[15] : r[479];
  assign _0053_ = sel_i[55] & ~(sel_i[54]);
  assign r_n[432] = _0053_ ? data_i[0] : r[448];
  assign r_n[433] = _0053_ ? data_i[1] : r[449];
  assign r_n[434] = _0053_ ? data_i[2] : r[450];
  assign r_n[435] = _0053_ ? data_i[3] : r[451];
  assign r_n[436] = _0053_ ? data_i[4] : r[452];
  assign r_n[437] = _0053_ ? data_i[5] : r[453];
  assign r_n[438] = _0053_ ? data_i[6] : r[454];
  assign r_n[439] = _0053_ ? data_i[7] : r[455];
  assign r_n[440] = _0053_ ? data_i[8] : r[456];
  assign r_n[441] = _0053_ ? data_i[9] : r[457];
  assign r_n[442] = _0053_ ? data_i[10] : r[458];
  assign r_n[443] = _0053_ ? data_i[11] : r[459];
  assign r_n[444] = _0053_ ? data_i[12] : r[460];
  assign r_n[445] = _0053_ ? data_i[13] : r[461];
  assign r_n[446] = _0053_ ? data_i[14] : r[462];
  assign r_n[447] = _0053_ ? data_i[15] : r[463];
  assign _0054_ = sel_i[53] & ~(sel_i[52]);
  assign r_n[416] = _0054_ ? data_i[0] : r[432];
  assign r_n[417] = _0054_ ? data_i[1] : r[433];
  assign r_n[418] = _0054_ ? data_i[2] : r[434];
  assign r_n[419] = _0054_ ? data_i[3] : r[435];
  assign r_n[420] = _0054_ ? data_i[4] : r[436];
  assign r_n[421] = _0054_ ? data_i[5] : r[437];
  assign r_n[422] = _0054_ ? data_i[6] : r[438];
  assign r_n[423] = _0054_ ? data_i[7] : r[439];
  assign r_n[424] = _0054_ ? data_i[8] : r[440];
  assign r_n[425] = _0054_ ? data_i[9] : r[441];
  assign r_n[426] = _0054_ ? data_i[10] : r[442];
  assign r_n[427] = _0054_ ? data_i[11] : r[443];
  assign r_n[428] = _0054_ ? data_i[12] : r[444];
  assign r_n[429] = _0054_ ? data_i[13] : r[445];
  assign r_n[430] = _0054_ ? data_i[14] : r[446];
  assign r_n[431] = _0054_ ? data_i[15] : r[447];
  assign _0055_ = sel_i[51] & ~(sel_i[50]);
  assign r_n[400] = _0055_ ? data_i[0] : r[416];
  assign r_n[401] = _0055_ ? data_i[1] : r[417];
  assign r_n[402] = _0055_ ? data_i[2] : r[418];
  assign r_n[403] = _0055_ ? data_i[3] : r[419];
  assign r_n[404] = _0055_ ? data_i[4] : r[420];
  assign r_n[405] = _0055_ ? data_i[5] : r[421];
  assign r_n[406] = _0055_ ? data_i[6] : r[422];
  assign r_n[407] = _0055_ ? data_i[7] : r[423];
  assign r_n[408] = _0055_ ? data_i[8] : r[424];
  assign r_n[409] = _0055_ ? data_i[9] : r[425];
  assign r_n[410] = _0055_ ? data_i[10] : r[426];
  assign r_n[411] = _0055_ ? data_i[11] : r[427];
  assign r_n[412] = _0055_ ? data_i[12] : r[428];
  assign r_n[413] = _0055_ ? data_i[13] : r[429];
  assign r_n[414] = _0055_ ? data_i[14] : r[430];
  assign r_n[415] = _0055_ ? data_i[15] : r[431];
  assign _0056_ = sel_i[49] & ~(sel_i[48]);
  assign r_n[384] = _0056_ ? data_i[0] : r[400];
  assign r_n[385] = _0056_ ? data_i[1] : r[401];
  assign r_n[386] = _0056_ ? data_i[2] : r[402];
  assign r_n[387] = _0056_ ? data_i[3] : r[403];
  assign r_n[388] = _0056_ ? data_i[4] : r[404];
  assign r_n[389] = _0056_ ? data_i[5] : r[405];
  assign r_n[390] = _0056_ ? data_i[6] : r[406];
  assign r_n[391] = _0056_ ? data_i[7] : r[407];
  assign r_n[392] = _0056_ ? data_i[8] : r[408];
  assign r_n[393] = _0056_ ? data_i[9] : r[409];
  assign r_n[394] = _0056_ ? data_i[10] : r[410];
  assign r_n[395] = _0056_ ? data_i[11] : r[411];
  assign r_n[396] = _0056_ ? data_i[12] : r[412];
  assign r_n[397] = _0056_ ? data_i[13] : r[413];
  assign r_n[398] = _0056_ ? data_i[14] : r[414];
  assign r_n[399] = _0056_ ? data_i[15] : r[415];
  assign _0057_ = sel_i[47] & ~(sel_i[46]);
  assign r_n[368] = _0057_ ? data_i[0] : r[384];
  assign r_n[369] = _0057_ ? data_i[1] : r[385];
  assign r_n[370] = _0057_ ? data_i[2] : r[386];
  assign r_n[371] = _0057_ ? data_i[3] : r[387];
  assign r_n[372] = _0057_ ? data_i[4] : r[388];
  assign r_n[373] = _0057_ ? data_i[5] : r[389];
  assign r_n[374] = _0057_ ? data_i[6] : r[390];
  assign r_n[375] = _0057_ ? data_i[7] : r[391];
  assign r_n[376] = _0057_ ? data_i[8] : r[392];
  assign r_n[377] = _0057_ ? data_i[9] : r[393];
  assign r_n[378] = _0057_ ? data_i[10] : r[394];
  assign r_n[379] = _0057_ ? data_i[11] : r[395];
  assign r_n[380] = _0057_ ? data_i[12] : r[396];
  assign r_n[381] = _0057_ ? data_i[13] : r[397];
  assign r_n[382] = _0057_ ? data_i[14] : r[398];
  assign r_n[383] = _0057_ ? data_i[15] : r[399];
  assign _0058_ = sel_i[45] & ~(sel_i[44]);
  assign r_n[352] = _0058_ ? data_i[0] : r[368];
  assign r_n[353] = _0058_ ? data_i[1] : r[369];
  assign r_n[354] = _0058_ ? data_i[2] : r[370];
  assign r_n[355] = _0058_ ? data_i[3] : r[371];
  assign r_n[356] = _0058_ ? data_i[4] : r[372];
  assign r_n[357] = _0058_ ? data_i[5] : r[373];
  assign r_n[358] = _0058_ ? data_i[6] : r[374];
  assign r_n[359] = _0058_ ? data_i[7] : r[375];
  assign r_n[360] = _0058_ ? data_i[8] : r[376];
  assign r_n[361] = _0058_ ? data_i[9] : r[377];
  assign r_n[362] = _0058_ ? data_i[10] : r[378];
  assign r_n[363] = _0058_ ? data_i[11] : r[379];
  assign r_n[364] = _0058_ ? data_i[12] : r[380];
  assign r_n[365] = _0058_ ? data_i[13] : r[381];
  assign r_n[366] = _0058_ ? data_i[14] : r[382];
  assign r_n[367] = _0058_ ? data_i[15] : r[383];
  assign _0059_ = sel_i[43] & ~(sel_i[42]);
  assign r_n[336] = _0059_ ? data_i[0] : r[352];
  assign r_n[337] = _0059_ ? data_i[1] : r[353];
  assign r_n[338] = _0059_ ? data_i[2] : r[354];
  assign r_n[339] = _0059_ ? data_i[3] : r[355];
  assign r_n[340] = _0059_ ? data_i[4] : r[356];
  assign r_n[341] = _0059_ ? data_i[5] : r[357];
  assign r_n[342] = _0059_ ? data_i[6] : r[358];
  assign r_n[343] = _0059_ ? data_i[7] : r[359];
  assign r_n[344] = _0059_ ? data_i[8] : r[360];
  assign r_n[345] = _0059_ ? data_i[9] : r[361];
  assign r_n[346] = _0059_ ? data_i[10] : r[362];
  assign r_n[347] = _0059_ ? data_i[11] : r[363];
  assign r_n[348] = _0059_ ? data_i[12] : r[364];
  assign r_n[349] = _0059_ ? data_i[13] : r[365];
  assign r_n[350] = _0059_ ? data_i[14] : r[366];
  assign r_n[351] = _0059_ ? data_i[15] : r[367];
  assign _0060_ = sel_i[41] & ~(sel_i[40]);
  assign r_n[320] = _0060_ ? data_i[0] : r[336];
  assign r_n[321] = _0060_ ? data_i[1] : r[337];
  assign r_n[322] = _0060_ ? data_i[2] : r[338];
  assign r_n[323] = _0060_ ? data_i[3] : r[339];
  assign r_n[324] = _0060_ ? data_i[4] : r[340];
  assign r_n[325] = _0060_ ? data_i[5] : r[341];
  assign r_n[326] = _0060_ ? data_i[6] : r[342];
  assign r_n[327] = _0060_ ? data_i[7] : r[343];
  assign r_n[328] = _0060_ ? data_i[8] : r[344];
  assign r_n[329] = _0060_ ? data_i[9] : r[345];
  assign r_n[330] = _0060_ ? data_i[10] : r[346];
  assign r_n[331] = _0060_ ? data_i[11] : r[347];
  assign r_n[332] = _0060_ ? data_i[12] : r[348];
  assign r_n[333] = _0060_ ? data_i[13] : r[349];
  assign r_n[334] = _0060_ ? data_i[14] : r[350];
  assign r_n[335] = _0060_ ? data_i[15] : r[351];
  assign _0061_ = sel_i[39] & ~(sel_i[38]);
  assign r_n[304] = _0061_ ? data_i[0] : r[320];
  assign r_n[305] = _0061_ ? data_i[1] : r[321];
  assign r_n[306] = _0061_ ? data_i[2] : r[322];
  assign r_n[307] = _0061_ ? data_i[3] : r[323];
  assign r_n[308] = _0061_ ? data_i[4] : r[324];
  assign r_n[309] = _0061_ ? data_i[5] : r[325];
  assign r_n[310] = _0061_ ? data_i[6] : r[326];
  assign r_n[311] = _0061_ ? data_i[7] : r[327];
  assign r_n[312] = _0061_ ? data_i[8] : r[328];
  assign r_n[313] = _0061_ ? data_i[9] : r[329];
  assign r_n[314] = _0061_ ? data_i[10] : r[330];
  assign r_n[315] = _0061_ ? data_i[11] : r[331];
  assign r_n[316] = _0061_ ? data_i[12] : r[332];
  assign r_n[317] = _0061_ ? data_i[13] : r[333];
  assign r_n[318] = _0061_ ? data_i[14] : r[334];
  assign r_n[319] = _0061_ ? data_i[15] : r[335];
  assign _0062_ = sel_i[37] & ~(sel_i[36]);
  assign r_n[288] = _0062_ ? data_i[0] : r[304];
  assign r_n[289] = _0062_ ? data_i[1] : r[305];
  assign r_n[290] = _0062_ ? data_i[2] : r[306];
  assign r_n[291] = _0062_ ? data_i[3] : r[307];
  assign r_n[292] = _0062_ ? data_i[4] : r[308];
  assign r_n[293] = _0062_ ? data_i[5] : r[309];
  assign r_n[294] = _0062_ ? data_i[6] : r[310];
  assign r_n[295] = _0062_ ? data_i[7] : r[311];
  assign r_n[296] = _0062_ ? data_i[8] : r[312];
  assign r_n[297] = _0062_ ? data_i[9] : r[313];
  assign r_n[298] = _0062_ ? data_i[10] : r[314];
  assign r_n[299] = _0062_ ? data_i[11] : r[315];
  assign r_n[300] = _0062_ ? data_i[12] : r[316];
  assign r_n[301] = _0062_ ? data_i[13] : r[317];
  assign r_n[302] = _0062_ ? data_i[14] : r[318];
  assign r_n[303] = _0062_ ? data_i[15] : r[319];
  assign _0063_ = sel_i[35] & ~(sel_i[34]);
  assign r_n[272] = _0063_ ? data_i[0] : r[288];
  assign r_n[273] = _0063_ ? data_i[1] : r[289];
  assign r_n[274] = _0063_ ? data_i[2] : r[290];
  assign r_n[275] = _0063_ ? data_i[3] : r[291];
  assign r_n[276] = _0063_ ? data_i[4] : r[292];
  assign r_n[277] = _0063_ ? data_i[5] : r[293];
  assign r_n[278] = _0063_ ? data_i[6] : r[294];
  assign r_n[279] = _0063_ ? data_i[7] : r[295];
  assign r_n[280] = _0063_ ? data_i[8] : r[296];
  assign r_n[281] = _0063_ ? data_i[9] : r[297];
  assign r_n[282] = _0063_ ? data_i[10] : r[298];
  assign r_n[283] = _0063_ ? data_i[11] : r[299];
  assign r_n[284] = _0063_ ? data_i[12] : r[300];
  assign r_n[285] = _0063_ ? data_i[13] : r[301];
  assign r_n[286] = _0063_ ? data_i[14] : r[302];
  assign r_n[287] = _0063_ ? data_i[15] : r[303];
  always @(posedge clk_i)
    if (_0000_) data_o[0] <= r_n[0];
  always @(posedge clk_i)
    if (_0000_) data_o[1] <= r_n[1];
  always @(posedge clk_i)
    if (_0000_) data_o[2] <= r_n[2];
  always @(posedge clk_i)
    if (_0000_) data_o[3] <= r_n[3];
  always @(posedge clk_i)
    if (_0000_) data_o[4] <= r_n[4];
  always @(posedge clk_i)
    if (_0000_) data_o[5] <= r_n[5];
  always @(posedge clk_i)
    if (_0000_) data_o[6] <= r_n[6];
  always @(posedge clk_i)
    if (_0000_) data_o[7] <= r_n[7];
  always @(posedge clk_i)
    if (_0000_) data_o[8] <= r_n[8];
  always @(posedge clk_i)
    if (_0000_) data_o[9] <= r_n[9];
  always @(posedge clk_i)
    if (_0000_) data_o[10] <= r_n[10];
  always @(posedge clk_i)
    if (_0000_) data_o[11] <= r_n[11];
  always @(posedge clk_i)
    if (_0000_) data_o[12] <= r_n[12];
  always @(posedge clk_i)
    if (_0000_) data_o[13] <= r_n[13];
  always @(posedge clk_i)
    if (_0000_) data_o[14] <= r_n[14];
  always @(posedge clk_i)
    if (_0000_) data_o[15] <= r_n[15];
  reg \r_reg[480] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[480]  <= r_n[480];
  assign r[480] = \r_reg[480] ;
  reg \r_reg[481] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[481]  <= r_n[481];
  assign r[481] = \r_reg[481] ;
  reg \r_reg[482] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[482]  <= r_n[482];
  assign r[482] = \r_reg[482] ;
  reg \r_reg[483] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[483]  <= r_n[483];
  assign r[483] = \r_reg[483] ;
  reg \r_reg[484] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[484]  <= r_n[484];
  assign r[484] = \r_reg[484] ;
  reg \r_reg[485] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[485]  <= r_n[485];
  assign r[485] = \r_reg[485] ;
  reg \r_reg[486] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[486]  <= r_n[486];
  assign r[486] = \r_reg[486] ;
  reg \r_reg[487] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[487]  <= r_n[487];
  assign r[487] = \r_reg[487] ;
  reg \r_reg[488] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[488]  <= r_n[488];
  assign r[488] = \r_reg[488] ;
  reg \r_reg[489] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[489]  <= r_n[489];
  assign r[489] = \r_reg[489] ;
  reg \r_reg[490] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[490]  <= r_n[490];
  assign r[490] = \r_reg[490] ;
  reg \r_reg[491] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[491]  <= r_n[491];
  assign r[491] = \r_reg[491] ;
  reg \r_reg[492] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[492]  <= r_n[492];
  assign r[492] = \r_reg[492] ;
  reg \r_reg[493] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[493]  <= r_n[493];
  assign r[493] = \r_reg[493] ;
  reg \r_reg[494] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[494]  <= r_n[494];
  assign r[494] = \r_reg[494] ;
  reg \r_reg[495] ;
  always @(posedge clk_i)
    if (_0030_) \r_reg[495]  <= r_n[495];
  assign r[495] = \r_reg[495] ;
  reg \r_reg[464] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[464]  <= r_n[464];
  assign r[464] = \r_reg[464] ;
  reg \r_reg[465] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[465]  <= r_n[465];
  assign r[465] = \r_reg[465] ;
  reg \r_reg[466] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[466]  <= r_n[466];
  assign r[466] = \r_reg[466] ;
  reg \r_reg[467] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[467]  <= r_n[467];
  assign r[467] = \r_reg[467] ;
  reg \r_reg[468] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[468]  <= r_n[468];
  assign r[468] = \r_reg[468] ;
  reg \r_reg[469] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[469]  <= r_n[469];
  assign r[469] = \r_reg[469] ;
  reg \r_reg[470] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[470]  <= r_n[470];
  assign r[470] = \r_reg[470] ;
  reg \r_reg[471] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[471]  <= r_n[471];
  assign r[471] = \r_reg[471] ;
  reg \r_reg[472] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[472]  <= r_n[472];
  assign r[472] = \r_reg[472] ;
  reg \r_reg[473] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[473]  <= r_n[473];
  assign r[473] = \r_reg[473] ;
  reg \r_reg[474] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[474]  <= r_n[474];
  assign r[474] = \r_reg[474] ;
  reg \r_reg[475] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[475]  <= r_n[475];
  assign r[475] = \r_reg[475] ;
  reg \r_reg[476] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[476]  <= r_n[476];
  assign r[476] = \r_reg[476] ;
  reg \r_reg[477] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[477]  <= r_n[477];
  assign r[477] = \r_reg[477] ;
  reg \r_reg[478] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[478]  <= r_n[478];
  assign r[478] = \r_reg[478] ;
  reg \r_reg[479] ;
  always @(posedge clk_i)
    if (_0029_) \r_reg[479]  <= r_n[479];
  assign r[479] = \r_reg[479] ;
  reg \r_reg[448] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[448]  <= r_n[448];
  assign r[448] = \r_reg[448] ;
  reg \r_reg[449] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[449]  <= r_n[449];
  assign r[449] = \r_reg[449] ;
  reg \r_reg[450] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[450]  <= r_n[450];
  assign r[450] = \r_reg[450] ;
  reg \r_reg[451] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[451]  <= r_n[451];
  assign r[451] = \r_reg[451] ;
  reg \r_reg[452] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[452]  <= r_n[452];
  assign r[452] = \r_reg[452] ;
  reg \r_reg[453] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[453]  <= r_n[453];
  assign r[453] = \r_reg[453] ;
  reg \r_reg[454] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[454]  <= r_n[454];
  assign r[454] = \r_reg[454] ;
  reg \r_reg[455] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[455]  <= r_n[455];
  assign r[455] = \r_reg[455] ;
  reg \r_reg[456] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[456]  <= r_n[456];
  assign r[456] = \r_reg[456] ;
  reg \r_reg[457] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[457]  <= r_n[457];
  assign r[457] = \r_reg[457] ;
  reg \r_reg[458] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[458]  <= r_n[458];
  assign r[458] = \r_reg[458] ;
  reg \r_reg[459] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[459]  <= r_n[459];
  assign r[459] = \r_reg[459] ;
  reg \r_reg[460] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[460]  <= r_n[460];
  assign r[460] = \r_reg[460] ;
  reg \r_reg[461] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[461]  <= r_n[461];
  assign r[461] = \r_reg[461] ;
  reg \r_reg[462] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[462]  <= r_n[462];
  assign r[462] = \r_reg[462] ;
  reg \r_reg[463] ;
  always @(posedge clk_i)
    if (_0028_) \r_reg[463]  <= r_n[463];
  assign r[463] = \r_reg[463] ;
  reg \r_reg[432] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[432]  <= r_n[432];
  assign r[432] = \r_reg[432] ;
  reg \r_reg[433] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[433]  <= r_n[433];
  assign r[433] = \r_reg[433] ;
  reg \r_reg[434] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[434]  <= r_n[434];
  assign r[434] = \r_reg[434] ;
  reg \r_reg[435] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[435]  <= r_n[435];
  assign r[435] = \r_reg[435] ;
  reg \r_reg[436] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[436]  <= r_n[436];
  assign r[436] = \r_reg[436] ;
  reg \r_reg[437] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[437]  <= r_n[437];
  assign r[437] = \r_reg[437] ;
  reg \r_reg[438] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[438]  <= r_n[438];
  assign r[438] = \r_reg[438] ;
  reg \r_reg[439] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[439]  <= r_n[439];
  assign r[439] = \r_reg[439] ;
  reg \r_reg[440] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[440]  <= r_n[440];
  assign r[440] = \r_reg[440] ;
  reg \r_reg[441] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[441]  <= r_n[441];
  assign r[441] = \r_reg[441] ;
  reg \r_reg[442] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[442]  <= r_n[442];
  assign r[442] = \r_reg[442] ;
  reg \r_reg[443] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[443]  <= r_n[443];
  assign r[443] = \r_reg[443] ;
  reg \r_reg[444] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[444]  <= r_n[444];
  assign r[444] = \r_reg[444] ;
  reg \r_reg[445] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[445]  <= r_n[445];
  assign r[445] = \r_reg[445] ;
  reg \r_reg[446] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[446]  <= r_n[446];
  assign r[446] = \r_reg[446] ;
  reg \r_reg[447] ;
  always @(posedge clk_i)
    if (_0027_) \r_reg[447]  <= r_n[447];
  assign r[447] = \r_reg[447] ;
  reg \r_reg[416] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[416]  <= r_n[416];
  assign r[416] = \r_reg[416] ;
  reg \r_reg[417] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[417]  <= r_n[417];
  assign r[417] = \r_reg[417] ;
  reg \r_reg[418] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[418]  <= r_n[418];
  assign r[418] = \r_reg[418] ;
  reg \r_reg[419] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[419]  <= r_n[419];
  assign r[419] = \r_reg[419] ;
  reg \r_reg[420] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[420]  <= r_n[420];
  assign r[420] = \r_reg[420] ;
  reg \r_reg[421] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[421]  <= r_n[421];
  assign r[421] = \r_reg[421] ;
  reg \r_reg[422] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[422]  <= r_n[422];
  assign r[422] = \r_reg[422] ;
  reg \r_reg[423] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[423]  <= r_n[423];
  assign r[423] = \r_reg[423] ;
  reg \r_reg[424] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[424]  <= r_n[424];
  assign r[424] = \r_reg[424] ;
  reg \r_reg[425] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[425]  <= r_n[425];
  assign r[425] = \r_reg[425] ;
  reg \r_reg[426] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[426]  <= r_n[426];
  assign r[426] = \r_reg[426] ;
  reg \r_reg[427] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[427]  <= r_n[427];
  assign r[427] = \r_reg[427] ;
  reg \r_reg[428] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[428]  <= r_n[428];
  assign r[428] = \r_reg[428] ;
  reg \r_reg[429] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[429]  <= r_n[429];
  assign r[429] = \r_reg[429] ;
  reg \r_reg[430] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[430]  <= r_n[430];
  assign r[430] = \r_reg[430] ;
  reg \r_reg[431] ;
  always @(posedge clk_i)
    if (_0026_) \r_reg[431]  <= r_n[431];
  assign r[431] = \r_reg[431] ;
  reg \r_reg[400] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[400]  <= r_n[400];
  assign r[400] = \r_reg[400] ;
  reg \r_reg[401] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[401]  <= r_n[401];
  assign r[401] = \r_reg[401] ;
  reg \r_reg[402] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[402]  <= r_n[402];
  assign r[402] = \r_reg[402] ;
  reg \r_reg[403] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[403]  <= r_n[403];
  assign r[403] = \r_reg[403] ;
  reg \r_reg[404] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[404]  <= r_n[404];
  assign r[404] = \r_reg[404] ;
  reg \r_reg[405] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[405]  <= r_n[405];
  assign r[405] = \r_reg[405] ;
  reg \r_reg[406] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[406]  <= r_n[406];
  assign r[406] = \r_reg[406] ;
  reg \r_reg[407] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[407]  <= r_n[407];
  assign r[407] = \r_reg[407] ;
  reg \r_reg[408] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[408]  <= r_n[408];
  assign r[408] = \r_reg[408] ;
  reg \r_reg[409] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[409]  <= r_n[409];
  assign r[409] = \r_reg[409] ;
  reg \r_reg[410] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[410]  <= r_n[410];
  assign r[410] = \r_reg[410] ;
  reg \r_reg[411] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[411]  <= r_n[411];
  assign r[411] = \r_reg[411] ;
  reg \r_reg[412] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[412]  <= r_n[412];
  assign r[412] = \r_reg[412] ;
  reg \r_reg[413] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[413]  <= r_n[413];
  assign r[413] = \r_reg[413] ;
  reg \r_reg[414] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[414]  <= r_n[414];
  assign r[414] = \r_reg[414] ;
  reg \r_reg[415] ;
  always @(posedge clk_i)
    if (_0025_) \r_reg[415]  <= r_n[415];
  assign r[415] = \r_reg[415] ;
  reg \r_reg[384] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[384]  <= r_n[384];
  assign r[384] = \r_reg[384] ;
  reg \r_reg[385] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[385]  <= r_n[385];
  assign r[385] = \r_reg[385] ;
  reg \r_reg[386] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[386]  <= r_n[386];
  assign r[386] = \r_reg[386] ;
  reg \r_reg[387] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[387]  <= r_n[387];
  assign r[387] = \r_reg[387] ;
  reg \r_reg[388] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[388]  <= r_n[388];
  assign r[388] = \r_reg[388] ;
  reg \r_reg[389] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[389]  <= r_n[389];
  assign r[389] = \r_reg[389] ;
  reg \r_reg[390] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[390]  <= r_n[390];
  assign r[390] = \r_reg[390] ;
  reg \r_reg[391] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[391]  <= r_n[391];
  assign r[391] = \r_reg[391] ;
  reg \r_reg[392] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[392]  <= r_n[392];
  assign r[392] = \r_reg[392] ;
  reg \r_reg[393] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[393]  <= r_n[393];
  assign r[393] = \r_reg[393] ;
  reg \r_reg[394] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[394]  <= r_n[394];
  assign r[394] = \r_reg[394] ;
  reg \r_reg[395] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[395]  <= r_n[395];
  assign r[395] = \r_reg[395] ;
  reg \r_reg[396] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[396]  <= r_n[396];
  assign r[396] = \r_reg[396] ;
  reg \r_reg[397] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[397]  <= r_n[397];
  assign r[397] = \r_reg[397] ;
  reg \r_reg[398] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[398]  <= r_n[398];
  assign r[398] = \r_reg[398] ;
  reg \r_reg[399] ;
  always @(posedge clk_i)
    if (_0024_) \r_reg[399]  <= r_n[399];
  assign r[399] = \r_reg[399] ;
  reg \r_reg[368] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[368]  <= r_n[368];
  assign r[368] = \r_reg[368] ;
  reg \r_reg[369] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[369]  <= r_n[369];
  assign r[369] = \r_reg[369] ;
  reg \r_reg[370] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[370]  <= r_n[370];
  assign r[370] = \r_reg[370] ;
  reg \r_reg[371] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[371]  <= r_n[371];
  assign r[371] = \r_reg[371] ;
  reg \r_reg[372] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[372]  <= r_n[372];
  assign r[372] = \r_reg[372] ;
  reg \r_reg[373] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[373]  <= r_n[373];
  assign r[373] = \r_reg[373] ;
  reg \r_reg[374] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[374]  <= r_n[374];
  assign r[374] = \r_reg[374] ;
  reg \r_reg[375] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[375]  <= r_n[375];
  assign r[375] = \r_reg[375] ;
  reg \r_reg[376] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[376]  <= r_n[376];
  assign r[376] = \r_reg[376] ;
  reg \r_reg[377] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[377]  <= r_n[377];
  assign r[377] = \r_reg[377] ;
  reg \r_reg[378] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[378]  <= r_n[378];
  assign r[378] = \r_reg[378] ;
  reg \r_reg[379] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[379]  <= r_n[379];
  assign r[379] = \r_reg[379] ;
  reg \r_reg[380] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[380]  <= r_n[380];
  assign r[380] = \r_reg[380] ;
  reg \r_reg[381] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[381]  <= r_n[381];
  assign r[381] = \r_reg[381] ;
  reg \r_reg[382] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[382]  <= r_n[382];
  assign r[382] = \r_reg[382] ;
  reg \r_reg[383] ;
  always @(posedge clk_i)
    if (_0023_) \r_reg[383]  <= r_n[383];
  assign r[383] = \r_reg[383] ;
  reg \r_reg[352] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[352]  <= r_n[352];
  assign r[352] = \r_reg[352] ;
  reg \r_reg[353] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[353]  <= r_n[353];
  assign r[353] = \r_reg[353] ;
  reg \r_reg[354] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[354]  <= r_n[354];
  assign r[354] = \r_reg[354] ;
  reg \r_reg[355] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[355]  <= r_n[355];
  assign r[355] = \r_reg[355] ;
  reg \r_reg[356] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[356]  <= r_n[356];
  assign r[356] = \r_reg[356] ;
  reg \r_reg[357] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[357]  <= r_n[357];
  assign r[357] = \r_reg[357] ;
  reg \r_reg[358] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[358]  <= r_n[358];
  assign r[358] = \r_reg[358] ;
  reg \r_reg[359] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[359]  <= r_n[359];
  assign r[359] = \r_reg[359] ;
  reg \r_reg[360] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[360]  <= r_n[360];
  assign r[360] = \r_reg[360] ;
  reg \r_reg[361] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[361]  <= r_n[361];
  assign r[361] = \r_reg[361] ;
  reg \r_reg[362] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[362]  <= r_n[362];
  assign r[362] = \r_reg[362] ;
  reg \r_reg[363] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[363]  <= r_n[363];
  assign r[363] = \r_reg[363] ;
  reg \r_reg[364] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[364]  <= r_n[364];
  assign r[364] = \r_reg[364] ;
  reg \r_reg[365] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[365]  <= r_n[365];
  assign r[365] = \r_reg[365] ;
  reg \r_reg[366] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[366]  <= r_n[366];
  assign r[366] = \r_reg[366] ;
  reg \r_reg[367] ;
  always @(posedge clk_i)
    if (_0022_) \r_reg[367]  <= r_n[367];
  assign r[367] = \r_reg[367] ;
  reg \r_reg[336] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[336]  <= r_n[336];
  assign r[336] = \r_reg[336] ;
  reg \r_reg[337] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[337]  <= r_n[337];
  assign r[337] = \r_reg[337] ;
  reg \r_reg[338] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[338]  <= r_n[338];
  assign r[338] = \r_reg[338] ;
  reg \r_reg[339] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[339]  <= r_n[339];
  assign r[339] = \r_reg[339] ;
  reg \r_reg[340] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[340]  <= r_n[340];
  assign r[340] = \r_reg[340] ;
  reg \r_reg[341] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[341]  <= r_n[341];
  assign r[341] = \r_reg[341] ;
  reg \r_reg[342] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[342]  <= r_n[342];
  assign r[342] = \r_reg[342] ;
  reg \r_reg[343] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[343]  <= r_n[343];
  assign r[343] = \r_reg[343] ;
  reg \r_reg[344] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[344]  <= r_n[344];
  assign r[344] = \r_reg[344] ;
  reg \r_reg[345] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[345]  <= r_n[345];
  assign r[345] = \r_reg[345] ;
  reg \r_reg[346] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[346]  <= r_n[346];
  assign r[346] = \r_reg[346] ;
  reg \r_reg[347] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[347]  <= r_n[347];
  assign r[347] = \r_reg[347] ;
  reg \r_reg[348] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[348]  <= r_n[348];
  assign r[348] = \r_reg[348] ;
  reg \r_reg[349] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[349]  <= r_n[349];
  assign r[349] = \r_reg[349] ;
  reg \r_reg[350] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[350]  <= r_n[350];
  assign r[350] = \r_reg[350] ;
  reg \r_reg[351] ;
  always @(posedge clk_i)
    if (_0021_) \r_reg[351]  <= r_n[351];
  assign r[351] = \r_reg[351] ;
  reg \r_reg[320] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[320]  <= r_n[320];
  assign r[320] = \r_reg[320] ;
  reg \r_reg[321] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[321]  <= r_n[321];
  assign r[321] = \r_reg[321] ;
  reg \r_reg[322] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[322]  <= r_n[322];
  assign r[322] = \r_reg[322] ;
  reg \r_reg[323] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[323]  <= r_n[323];
  assign r[323] = \r_reg[323] ;
  reg \r_reg[324] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[324]  <= r_n[324];
  assign r[324] = \r_reg[324] ;
  reg \r_reg[325] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[325]  <= r_n[325];
  assign r[325] = \r_reg[325] ;
  reg \r_reg[326] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[326]  <= r_n[326];
  assign r[326] = \r_reg[326] ;
  reg \r_reg[327] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[327]  <= r_n[327];
  assign r[327] = \r_reg[327] ;
  reg \r_reg[328] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[328]  <= r_n[328];
  assign r[328] = \r_reg[328] ;
  reg \r_reg[329] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[329]  <= r_n[329];
  assign r[329] = \r_reg[329] ;
  reg \r_reg[330] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[330]  <= r_n[330];
  assign r[330] = \r_reg[330] ;
  reg \r_reg[331] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[331]  <= r_n[331];
  assign r[331] = \r_reg[331] ;
  reg \r_reg[332] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[332]  <= r_n[332];
  assign r[332] = \r_reg[332] ;
  reg \r_reg[333] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[333]  <= r_n[333];
  assign r[333] = \r_reg[333] ;
  reg \r_reg[334] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[334]  <= r_n[334];
  assign r[334] = \r_reg[334] ;
  reg \r_reg[335] ;
  always @(posedge clk_i)
    if (_0020_) \r_reg[335]  <= r_n[335];
  assign r[335] = \r_reg[335] ;
  reg \r_reg[304] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[304]  <= r_n[304];
  assign r[304] = \r_reg[304] ;
  reg \r_reg[305] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[305]  <= r_n[305];
  assign r[305] = \r_reg[305] ;
  reg \r_reg[306] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[306]  <= r_n[306];
  assign r[306] = \r_reg[306] ;
  reg \r_reg[307] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[307]  <= r_n[307];
  assign r[307] = \r_reg[307] ;
  reg \r_reg[308] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[308]  <= r_n[308];
  assign r[308] = \r_reg[308] ;
  reg \r_reg[309] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[309]  <= r_n[309];
  assign r[309] = \r_reg[309] ;
  reg \r_reg[310] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[310]  <= r_n[310];
  assign r[310] = \r_reg[310] ;
  reg \r_reg[311] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[311]  <= r_n[311];
  assign r[311] = \r_reg[311] ;
  reg \r_reg[312] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[312]  <= r_n[312];
  assign r[312] = \r_reg[312] ;
  reg \r_reg[313] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[313]  <= r_n[313];
  assign r[313] = \r_reg[313] ;
  reg \r_reg[314] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[314]  <= r_n[314];
  assign r[314] = \r_reg[314] ;
  reg \r_reg[315] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[315]  <= r_n[315];
  assign r[315] = \r_reg[315] ;
  reg \r_reg[316] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[316]  <= r_n[316];
  assign r[316] = \r_reg[316] ;
  reg \r_reg[317] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[317]  <= r_n[317];
  assign r[317] = \r_reg[317] ;
  reg \r_reg[318] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[318]  <= r_n[318];
  assign r[318] = \r_reg[318] ;
  reg \r_reg[319] ;
  always @(posedge clk_i)
    if (_0019_) \r_reg[319]  <= r_n[319];
  assign r[319] = \r_reg[319] ;
  reg \r_reg[288] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[288]  <= r_n[288];
  assign r[288] = \r_reg[288] ;
  reg \r_reg[289] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[289]  <= r_n[289];
  assign r[289] = \r_reg[289] ;
  reg \r_reg[290] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[290]  <= r_n[290];
  assign r[290] = \r_reg[290] ;
  reg \r_reg[291] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[291]  <= r_n[291];
  assign r[291] = \r_reg[291] ;
  reg \r_reg[292] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[292]  <= r_n[292];
  assign r[292] = \r_reg[292] ;
  reg \r_reg[293] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[293]  <= r_n[293];
  assign r[293] = \r_reg[293] ;
  reg \r_reg[294] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[294]  <= r_n[294];
  assign r[294] = \r_reg[294] ;
  reg \r_reg[295] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[295]  <= r_n[295];
  assign r[295] = \r_reg[295] ;
  reg \r_reg[296] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[296]  <= r_n[296];
  assign r[296] = \r_reg[296] ;
  reg \r_reg[297] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[297]  <= r_n[297];
  assign r[297] = \r_reg[297] ;
  reg \r_reg[298] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[298]  <= r_n[298];
  assign r[298] = \r_reg[298] ;
  reg \r_reg[299] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[299]  <= r_n[299];
  assign r[299] = \r_reg[299] ;
  reg \r_reg[300] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[300]  <= r_n[300];
  assign r[300] = \r_reg[300] ;
  reg \r_reg[301] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[301]  <= r_n[301];
  assign r[301] = \r_reg[301] ;
  reg \r_reg[302] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[302]  <= r_n[302];
  assign r[302] = \r_reg[302] ;
  reg \r_reg[303] ;
  always @(posedge clk_i)
    if (_0018_) \r_reg[303]  <= r_n[303];
  assign r[303] = \r_reg[303] ;
  reg \r_reg[272] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[272]  <= r_n[272];
  assign r[272] = \r_reg[272] ;
  reg \r_reg[273] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[273]  <= r_n[273];
  assign r[273] = \r_reg[273] ;
  reg \r_reg[274] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[274]  <= r_n[274];
  assign r[274] = \r_reg[274] ;
  reg \r_reg[275] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[275]  <= r_n[275];
  assign r[275] = \r_reg[275] ;
  reg \r_reg[276] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[276]  <= r_n[276];
  assign r[276] = \r_reg[276] ;
  reg \r_reg[277] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[277]  <= r_n[277];
  assign r[277] = \r_reg[277] ;
  reg \r_reg[278] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[278]  <= r_n[278];
  assign r[278] = \r_reg[278] ;
  reg \r_reg[279] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[279]  <= r_n[279];
  assign r[279] = \r_reg[279] ;
  reg \r_reg[280] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[280]  <= r_n[280];
  assign r[280] = \r_reg[280] ;
  reg \r_reg[281] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[281]  <= r_n[281];
  assign r[281] = \r_reg[281] ;
  reg \r_reg[282] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[282]  <= r_n[282];
  assign r[282] = \r_reg[282] ;
  reg \r_reg[283] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[283]  <= r_n[283];
  assign r[283] = \r_reg[283] ;
  reg \r_reg[284] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[284]  <= r_n[284];
  assign r[284] = \r_reg[284] ;
  reg \r_reg[285] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[285]  <= r_n[285];
  assign r[285] = \r_reg[285] ;
  reg \r_reg[286] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[286]  <= r_n[286];
  assign r[286] = \r_reg[286] ;
  reg \r_reg[287] ;
  always @(posedge clk_i)
    if (_0017_) \r_reg[287]  <= r_n[287];
  assign r[287] = \r_reg[287] ;
  reg \r_reg[256] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[256]  <= r_n[256];
  assign r[256] = \r_reg[256] ;
  reg \r_reg[257] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[257]  <= r_n[257];
  assign r[257] = \r_reg[257] ;
  reg \r_reg[258] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[258]  <= r_n[258];
  assign r[258] = \r_reg[258] ;
  reg \r_reg[259] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[259]  <= r_n[259];
  assign r[259] = \r_reg[259] ;
  reg \r_reg[260] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[260]  <= r_n[260];
  assign r[260] = \r_reg[260] ;
  reg \r_reg[261] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[261]  <= r_n[261];
  assign r[261] = \r_reg[261] ;
  reg \r_reg[262] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[262]  <= r_n[262];
  assign r[262] = \r_reg[262] ;
  reg \r_reg[263] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[263]  <= r_n[263];
  assign r[263] = \r_reg[263] ;
  reg \r_reg[264] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[264]  <= r_n[264];
  assign r[264] = \r_reg[264] ;
  reg \r_reg[265] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[265]  <= r_n[265];
  assign r[265] = \r_reg[265] ;
  reg \r_reg[266] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[266]  <= r_n[266];
  assign r[266] = \r_reg[266] ;
  reg \r_reg[267] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[267]  <= r_n[267];
  assign r[267] = \r_reg[267] ;
  reg \r_reg[268] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[268]  <= r_n[268];
  assign r[268] = \r_reg[268] ;
  reg \r_reg[269] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[269]  <= r_n[269];
  assign r[269] = \r_reg[269] ;
  reg \r_reg[270] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[270]  <= r_n[270];
  assign r[270] = \r_reg[270] ;
  reg \r_reg[271] ;
  always @(posedge clk_i)
    if (_0016_) \r_reg[271]  <= r_n[271];
  assign r[271] = \r_reg[271] ;
  reg \r_reg[240] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[240]  <= r_n[240];
  assign r[240] = \r_reg[240] ;
  reg \r_reg[241] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[241]  <= r_n[241];
  assign r[241] = \r_reg[241] ;
  reg \r_reg[242] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[242]  <= r_n[242];
  assign r[242] = \r_reg[242] ;
  reg \r_reg[243] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[243]  <= r_n[243];
  assign r[243] = \r_reg[243] ;
  reg \r_reg[244] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[244]  <= r_n[244];
  assign r[244] = \r_reg[244] ;
  reg \r_reg[245] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[245]  <= r_n[245];
  assign r[245] = \r_reg[245] ;
  reg \r_reg[246] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[246]  <= r_n[246];
  assign r[246] = \r_reg[246] ;
  reg \r_reg[247] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[247]  <= r_n[247];
  assign r[247] = \r_reg[247] ;
  reg \r_reg[248] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[248]  <= r_n[248];
  assign r[248] = \r_reg[248] ;
  reg \r_reg[249] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[249]  <= r_n[249];
  assign r[249] = \r_reg[249] ;
  reg \r_reg[250] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[250]  <= r_n[250];
  assign r[250] = \r_reg[250] ;
  reg \r_reg[251] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[251]  <= r_n[251];
  assign r[251] = \r_reg[251] ;
  reg \r_reg[252] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[252]  <= r_n[252];
  assign r[252] = \r_reg[252] ;
  reg \r_reg[253] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[253]  <= r_n[253];
  assign r[253] = \r_reg[253] ;
  reg \r_reg[254] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[254]  <= r_n[254];
  assign r[254] = \r_reg[254] ;
  reg \r_reg[255] ;
  always @(posedge clk_i)
    if (_0015_) \r_reg[255]  <= r_n[255];
  assign r[255] = \r_reg[255] ;
  reg \r_reg[224] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[224]  <= r_n[224];
  assign r[224] = \r_reg[224] ;
  reg \r_reg[225] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[225]  <= r_n[225];
  assign r[225] = \r_reg[225] ;
  reg \r_reg[226] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[226]  <= r_n[226];
  assign r[226] = \r_reg[226] ;
  reg \r_reg[227] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[227]  <= r_n[227];
  assign r[227] = \r_reg[227] ;
  reg \r_reg[228] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[228]  <= r_n[228];
  assign r[228] = \r_reg[228] ;
  reg \r_reg[229] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[229]  <= r_n[229];
  assign r[229] = \r_reg[229] ;
  reg \r_reg[230] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[230]  <= r_n[230];
  assign r[230] = \r_reg[230] ;
  reg \r_reg[231] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[231]  <= r_n[231];
  assign r[231] = \r_reg[231] ;
  reg \r_reg[232] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[232]  <= r_n[232];
  assign r[232] = \r_reg[232] ;
  reg \r_reg[233] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[233]  <= r_n[233];
  assign r[233] = \r_reg[233] ;
  reg \r_reg[234] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[234]  <= r_n[234];
  assign r[234] = \r_reg[234] ;
  reg \r_reg[235] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[235]  <= r_n[235];
  assign r[235] = \r_reg[235] ;
  reg \r_reg[236] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[236]  <= r_n[236];
  assign r[236] = \r_reg[236] ;
  reg \r_reg[237] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[237]  <= r_n[237];
  assign r[237] = \r_reg[237] ;
  reg \r_reg[238] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[238]  <= r_n[238];
  assign r[238] = \r_reg[238] ;
  reg \r_reg[239] ;
  always @(posedge clk_i)
    if (_0014_) \r_reg[239]  <= r_n[239];
  assign r[239] = \r_reg[239] ;
  reg \r_reg[208] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[208]  <= r_n[208];
  assign r[208] = \r_reg[208] ;
  reg \r_reg[209] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[209]  <= r_n[209];
  assign r[209] = \r_reg[209] ;
  reg \r_reg[210] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[210]  <= r_n[210];
  assign r[210] = \r_reg[210] ;
  reg \r_reg[211] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[211]  <= r_n[211];
  assign r[211] = \r_reg[211] ;
  reg \r_reg[212] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[212]  <= r_n[212];
  assign r[212] = \r_reg[212] ;
  reg \r_reg[213] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[213]  <= r_n[213];
  assign r[213] = \r_reg[213] ;
  reg \r_reg[214] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[214]  <= r_n[214];
  assign r[214] = \r_reg[214] ;
  reg \r_reg[215] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[215]  <= r_n[215];
  assign r[215] = \r_reg[215] ;
  reg \r_reg[216] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[216]  <= r_n[216];
  assign r[216] = \r_reg[216] ;
  reg \r_reg[217] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[217]  <= r_n[217];
  assign r[217] = \r_reg[217] ;
  reg \r_reg[218] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[218]  <= r_n[218];
  assign r[218] = \r_reg[218] ;
  reg \r_reg[219] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[219]  <= r_n[219];
  assign r[219] = \r_reg[219] ;
  reg \r_reg[220] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[220]  <= r_n[220];
  assign r[220] = \r_reg[220] ;
  reg \r_reg[221] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[221]  <= r_n[221];
  assign r[221] = \r_reg[221] ;
  reg \r_reg[222] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[222]  <= r_n[222];
  assign r[222] = \r_reg[222] ;
  reg \r_reg[223] ;
  always @(posedge clk_i)
    if (_0013_) \r_reg[223]  <= r_n[223];
  assign r[223] = \r_reg[223] ;
  reg \r_reg[192] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[192]  <= r_n[192];
  assign r[192] = \r_reg[192] ;
  reg \r_reg[193] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[193]  <= r_n[193];
  assign r[193] = \r_reg[193] ;
  reg \r_reg[194] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[194]  <= r_n[194];
  assign r[194] = \r_reg[194] ;
  reg \r_reg[195] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[195]  <= r_n[195];
  assign r[195] = \r_reg[195] ;
  reg \r_reg[196] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[196]  <= r_n[196];
  assign r[196] = \r_reg[196] ;
  reg \r_reg[197] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[197]  <= r_n[197];
  assign r[197] = \r_reg[197] ;
  reg \r_reg[198] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[198]  <= r_n[198];
  assign r[198] = \r_reg[198] ;
  reg \r_reg[199] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[199]  <= r_n[199];
  assign r[199] = \r_reg[199] ;
  reg \r_reg[200] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[200]  <= r_n[200];
  assign r[200] = \r_reg[200] ;
  reg \r_reg[201] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[201]  <= r_n[201];
  assign r[201] = \r_reg[201] ;
  reg \r_reg[202] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[202]  <= r_n[202];
  assign r[202] = \r_reg[202] ;
  reg \r_reg[203] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[203]  <= r_n[203];
  assign r[203] = \r_reg[203] ;
  reg \r_reg[204] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[204]  <= r_n[204];
  assign r[204] = \r_reg[204] ;
  reg \r_reg[205] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[205]  <= r_n[205];
  assign r[205] = \r_reg[205] ;
  reg \r_reg[206] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[206]  <= r_n[206];
  assign r[206] = \r_reg[206] ;
  reg \r_reg[207] ;
  always @(posedge clk_i)
    if (_0012_) \r_reg[207]  <= r_n[207];
  assign r[207] = \r_reg[207] ;
  reg \r_reg[176] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[176]  <= r_n[176];
  assign r[176] = \r_reg[176] ;
  reg \r_reg[177] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[177]  <= r_n[177];
  assign r[177] = \r_reg[177] ;
  reg \r_reg[178] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[178]  <= r_n[178];
  assign r[178] = \r_reg[178] ;
  reg \r_reg[179] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[179]  <= r_n[179];
  assign r[179] = \r_reg[179] ;
  reg \r_reg[180] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[180]  <= r_n[180];
  assign r[180] = \r_reg[180] ;
  reg \r_reg[181] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[181]  <= r_n[181];
  assign r[181] = \r_reg[181] ;
  reg \r_reg[182] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[182]  <= r_n[182];
  assign r[182] = \r_reg[182] ;
  reg \r_reg[183] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[183]  <= r_n[183];
  assign r[183] = \r_reg[183] ;
  reg \r_reg[184] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[184]  <= r_n[184];
  assign r[184] = \r_reg[184] ;
  reg \r_reg[185] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[185]  <= r_n[185];
  assign r[185] = \r_reg[185] ;
  reg \r_reg[186] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[186]  <= r_n[186];
  assign r[186] = \r_reg[186] ;
  reg \r_reg[187] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[187]  <= r_n[187];
  assign r[187] = \r_reg[187] ;
  reg \r_reg[188] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[188]  <= r_n[188];
  assign r[188] = \r_reg[188] ;
  reg \r_reg[189] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[189]  <= r_n[189];
  assign r[189] = \r_reg[189] ;
  reg \r_reg[190] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[190]  <= r_n[190];
  assign r[190] = \r_reg[190] ;
  reg \r_reg[191] ;
  always @(posedge clk_i)
    if (_0011_) \r_reg[191]  <= r_n[191];
  assign r[191] = \r_reg[191] ;
  reg \r_reg[160] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[160]  <= r_n[160];
  assign r[160] = \r_reg[160] ;
  reg \r_reg[161] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[161]  <= r_n[161];
  assign r[161] = \r_reg[161] ;
  reg \r_reg[162] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[162]  <= r_n[162];
  assign r[162] = \r_reg[162] ;
  reg \r_reg[163] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[163]  <= r_n[163];
  assign r[163] = \r_reg[163] ;
  reg \r_reg[164] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[164]  <= r_n[164];
  assign r[164] = \r_reg[164] ;
  reg \r_reg[165] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[165]  <= r_n[165];
  assign r[165] = \r_reg[165] ;
  reg \r_reg[166] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[166]  <= r_n[166];
  assign r[166] = \r_reg[166] ;
  reg \r_reg[167] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[167]  <= r_n[167];
  assign r[167] = \r_reg[167] ;
  reg \r_reg[168] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[168]  <= r_n[168];
  assign r[168] = \r_reg[168] ;
  reg \r_reg[169] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[169]  <= r_n[169];
  assign r[169] = \r_reg[169] ;
  reg \r_reg[170] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[170]  <= r_n[170];
  assign r[170] = \r_reg[170] ;
  reg \r_reg[171] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[171]  <= r_n[171];
  assign r[171] = \r_reg[171] ;
  reg \r_reg[172] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[172]  <= r_n[172];
  assign r[172] = \r_reg[172] ;
  reg \r_reg[173] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[173]  <= r_n[173];
  assign r[173] = \r_reg[173] ;
  reg \r_reg[174] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[174]  <= r_n[174];
  assign r[174] = \r_reg[174] ;
  reg \r_reg[175] ;
  always @(posedge clk_i)
    if (_0010_) \r_reg[175]  <= r_n[175];
  assign r[175] = \r_reg[175] ;
  reg \r_reg[144] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[144]  <= r_n[144];
  assign r[144] = \r_reg[144] ;
  reg \r_reg[145] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[145]  <= r_n[145];
  assign r[145] = \r_reg[145] ;
  reg \r_reg[146] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[146]  <= r_n[146];
  assign r[146] = \r_reg[146] ;
  reg \r_reg[147] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[147]  <= r_n[147];
  assign r[147] = \r_reg[147] ;
  reg \r_reg[148] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[148]  <= r_n[148];
  assign r[148] = \r_reg[148] ;
  reg \r_reg[149] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[149]  <= r_n[149];
  assign r[149] = \r_reg[149] ;
  reg \r_reg[150] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[150]  <= r_n[150];
  assign r[150] = \r_reg[150] ;
  reg \r_reg[151] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[151]  <= r_n[151];
  assign r[151] = \r_reg[151] ;
  reg \r_reg[152] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[152]  <= r_n[152];
  assign r[152] = \r_reg[152] ;
  reg \r_reg[153] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[153]  <= r_n[153];
  assign r[153] = \r_reg[153] ;
  reg \r_reg[154] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[154]  <= r_n[154];
  assign r[154] = \r_reg[154] ;
  reg \r_reg[155] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[155]  <= r_n[155];
  assign r[155] = \r_reg[155] ;
  reg \r_reg[156] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[156]  <= r_n[156];
  assign r[156] = \r_reg[156] ;
  reg \r_reg[157] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[157]  <= r_n[157];
  assign r[157] = \r_reg[157] ;
  reg \r_reg[158] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[158]  <= r_n[158];
  assign r[158] = \r_reg[158] ;
  reg \r_reg[159] ;
  always @(posedge clk_i)
    if (_0009_) \r_reg[159]  <= r_n[159];
  assign r[159] = \r_reg[159] ;
  reg \r_reg[128] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[128]  <= r_n[128];
  assign r[128] = \r_reg[128] ;
  reg \r_reg[129] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[129]  <= r_n[129];
  assign r[129] = \r_reg[129] ;
  reg \r_reg[130] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[130]  <= r_n[130];
  assign r[130] = \r_reg[130] ;
  reg \r_reg[131] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[131]  <= r_n[131];
  assign r[131] = \r_reg[131] ;
  reg \r_reg[132] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[132]  <= r_n[132];
  assign r[132] = \r_reg[132] ;
  reg \r_reg[133] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[133]  <= r_n[133];
  assign r[133] = \r_reg[133] ;
  reg \r_reg[134] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[134]  <= r_n[134];
  assign r[134] = \r_reg[134] ;
  reg \r_reg[135] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[135]  <= r_n[135];
  assign r[135] = \r_reg[135] ;
  reg \r_reg[136] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[136]  <= r_n[136];
  assign r[136] = \r_reg[136] ;
  reg \r_reg[137] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[137]  <= r_n[137];
  assign r[137] = \r_reg[137] ;
  reg \r_reg[138] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[138]  <= r_n[138];
  assign r[138] = \r_reg[138] ;
  reg \r_reg[139] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[139]  <= r_n[139];
  assign r[139] = \r_reg[139] ;
  reg \r_reg[140] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[140]  <= r_n[140];
  assign r[140] = \r_reg[140] ;
  reg \r_reg[141] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[141]  <= r_n[141];
  assign r[141] = \r_reg[141] ;
  reg \r_reg[142] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[142]  <= r_n[142];
  assign r[142] = \r_reg[142] ;
  reg \r_reg[143] ;
  always @(posedge clk_i)
    if (_0008_) \r_reg[143]  <= r_n[143];
  assign r[143] = \r_reg[143] ;
  reg \r_reg[112] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[112]  <= r_n[112];
  assign r[112] = \r_reg[112] ;
  reg \r_reg[113] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[113]  <= r_n[113];
  assign r[113] = \r_reg[113] ;
  reg \r_reg[114] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[114]  <= r_n[114];
  assign r[114] = \r_reg[114] ;
  reg \r_reg[115] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[115]  <= r_n[115];
  assign r[115] = \r_reg[115] ;
  reg \r_reg[116] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[116]  <= r_n[116];
  assign r[116] = \r_reg[116] ;
  reg \r_reg[117] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[117]  <= r_n[117];
  assign r[117] = \r_reg[117] ;
  reg \r_reg[118] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[118]  <= r_n[118];
  assign r[118] = \r_reg[118] ;
  reg \r_reg[119] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[119]  <= r_n[119];
  assign r[119] = \r_reg[119] ;
  reg \r_reg[120] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[120]  <= r_n[120];
  assign r[120] = \r_reg[120] ;
  reg \r_reg[121] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[121]  <= r_n[121];
  assign r[121] = \r_reg[121] ;
  reg \r_reg[122] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[122]  <= r_n[122];
  assign r[122] = \r_reg[122] ;
  reg \r_reg[123] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[123]  <= r_n[123];
  assign r[123] = \r_reg[123] ;
  reg \r_reg[124] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[124]  <= r_n[124];
  assign r[124] = \r_reg[124] ;
  reg \r_reg[125] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[125]  <= r_n[125];
  assign r[125] = \r_reg[125] ;
  reg \r_reg[126] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[126]  <= r_n[126];
  assign r[126] = \r_reg[126] ;
  reg \r_reg[127] ;
  always @(posedge clk_i)
    if (_0007_) \r_reg[127]  <= r_n[127];
  assign r[127] = \r_reg[127] ;
  reg \r_reg[96] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[96]  <= r_n[96];
  assign r[96] = \r_reg[96] ;
  reg \r_reg[97] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[97]  <= r_n[97];
  assign r[97] = \r_reg[97] ;
  reg \r_reg[98] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[98]  <= r_n[98];
  assign r[98] = \r_reg[98] ;
  reg \r_reg[99] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[99]  <= r_n[99];
  assign r[99] = \r_reg[99] ;
  reg \r_reg[100] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[100]  <= r_n[100];
  assign r[100] = \r_reg[100] ;
  reg \r_reg[101] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[101]  <= r_n[101];
  assign r[101] = \r_reg[101] ;
  reg \r_reg[102] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[102]  <= r_n[102];
  assign r[102] = \r_reg[102] ;
  reg \r_reg[103] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[103]  <= r_n[103];
  assign r[103] = \r_reg[103] ;
  reg \r_reg[104] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[104]  <= r_n[104];
  assign r[104] = \r_reg[104] ;
  reg \r_reg[105] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[105]  <= r_n[105];
  assign r[105] = \r_reg[105] ;
  reg \r_reg[106] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[106]  <= r_n[106];
  assign r[106] = \r_reg[106] ;
  reg \r_reg[107] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[107]  <= r_n[107];
  assign r[107] = \r_reg[107] ;
  reg \r_reg[108] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[108]  <= r_n[108];
  assign r[108] = \r_reg[108] ;
  reg \r_reg[109] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[109]  <= r_n[109];
  assign r[109] = \r_reg[109] ;
  reg \r_reg[110] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[110]  <= r_n[110];
  assign r[110] = \r_reg[110] ;
  reg \r_reg[111] ;
  always @(posedge clk_i)
    if (_0006_) \r_reg[111]  <= r_n[111];
  assign r[111] = \r_reg[111] ;
  reg \r_reg[80] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[80]  <= r_n[80];
  assign r[80] = \r_reg[80] ;
  reg \r_reg[81] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[81]  <= r_n[81];
  assign r[81] = \r_reg[81] ;
  reg \r_reg[82] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[82]  <= r_n[82];
  assign r[82] = \r_reg[82] ;
  reg \r_reg[83] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[83]  <= r_n[83];
  assign r[83] = \r_reg[83] ;
  reg \r_reg[84] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[84]  <= r_n[84];
  assign r[84] = \r_reg[84] ;
  reg \r_reg[85] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[85]  <= r_n[85];
  assign r[85] = \r_reg[85] ;
  reg \r_reg[86] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[86]  <= r_n[86];
  assign r[86] = \r_reg[86] ;
  reg \r_reg[87] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[87]  <= r_n[87];
  assign r[87] = \r_reg[87] ;
  reg \r_reg[88] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[88]  <= r_n[88];
  assign r[88] = \r_reg[88] ;
  reg \r_reg[89] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[89]  <= r_n[89];
  assign r[89] = \r_reg[89] ;
  reg \r_reg[90] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[90]  <= r_n[90];
  assign r[90] = \r_reg[90] ;
  reg \r_reg[91] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[91]  <= r_n[91];
  assign r[91] = \r_reg[91] ;
  reg \r_reg[92] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[92]  <= r_n[92];
  assign r[92] = \r_reg[92] ;
  reg \r_reg[93] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[93]  <= r_n[93];
  assign r[93] = \r_reg[93] ;
  reg \r_reg[94] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[94]  <= r_n[94];
  assign r[94] = \r_reg[94] ;
  reg \r_reg[95] ;
  always @(posedge clk_i)
    if (_0005_) \r_reg[95]  <= r_n[95];
  assign r[95] = \r_reg[95] ;
  reg \r_reg[64] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[64]  <= r_n[64];
  assign r[64] = \r_reg[64] ;
  reg \r_reg[65] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[65]  <= r_n[65];
  assign r[65] = \r_reg[65] ;
  reg \r_reg[66] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[66]  <= r_n[66];
  assign r[66] = \r_reg[66] ;
  reg \r_reg[67] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[67]  <= r_n[67];
  assign r[67] = \r_reg[67] ;
  reg \r_reg[68] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[68]  <= r_n[68];
  assign r[68] = \r_reg[68] ;
  reg \r_reg[69] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[69]  <= r_n[69];
  assign r[69] = \r_reg[69] ;
  reg \r_reg[70] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[70]  <= r_n[70];
  assign r[70] = \r_reg[70] ;
  reg \r_reg[71] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[71]  <= r_n[71];
  assign r[71] = \r_reg[71] ;
  reg \r_reg[72] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[72]  <= r_n[72];
  assign r[72] = \r_reg[72] ;
  reg \r_reg[73] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[73]  <= r_n[73];
  assign r[73] = \r_reg[73] ;
  reg \r_reg[74] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[74]  <= r_n[74];
  assign r[74] = \r_reg[74] ;
  reg \r_reg[75] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[75]  <= r_n[75];
  assign r[75] = \r_reg[75] ;
  reg \r_reg[76] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[76]  <= r_n[76];
  assign r[76] = \r_reg[76] ;
  reg \r_reg[77] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[77]  <= r_n[77];
  assign r[77] = \r_reg[77] ;
  reg \r_reg[78] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[78]  <= r_n[78];
  assign r[78] = \r_reg[78] ;
  reg \r_reg[79] ;
  always @(posedge clk_i)
    if (_0004_) \r_reg[79]  <= r_n[79];
  assign r[79] = \r_reg[79] ;
  reg \r_reg[48] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[48]  <= r_n[48];
  assign r[48] = \r_reg[48] ;
  reg \r_reg[49] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[49]  <= r_n[49];
  assign r[49] = \r_reg[49] ;
  reg \r_reg[50] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[50]  <= r_n[50];
  assign r[50] = \r_reg[50] ;
  reg \r_reg[51] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[51]  <= r_n[51];
  assign r[51] = \r_reg[51] ;
  reg \r_reg[52] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[52]  <= r_n[52];
  assign r[52] = \r_reg[52] ;
  reg \r_reg[53] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[53]  <= r_n[53];
  assign r[53] = \r_reg[53] ;
  reg \r_reg[54] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[54]  <= r_n[54];
  assign r[54] = \r_reg[54] ;
  reg \r_reg[55] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[55]  <= r_n[55];
  assign r[55] = \r_reg[55] ;
  reg \r_reg[56] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[56]  <= r_n[56];
  assign r[56] = \r_reg[56] ;
  reg \r_reg[57] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[57]  <= r_n[57];
  assign r[57] = \r_reg[57] ;
  reg \r_reg[58] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[58]  <= r_n[58];
  assign r[58] = \r_reg[58] ;
  reg \r_reg[59] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[59]  <= r_n[59];
  assign r[59] = \r_reg[59] ;
  reg \r_reg[60] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[60]  <= r_n[60];
  assign r[60] = \r_reg[60] ;
  reg \r_reg[61] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[61]  <= r_n[61];
  assign r[61] = \r_reg[61] ;
  reg \r_reg[62] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[62]  <= r_n[62];
  assign r[62] = \r_reg[62] ;
  reg \r_reg[63] ;
  always @(posedge clk_i)
    if (_0003_) \r_reg[63]  <= r_n[63];
  assign r[63] = \r_reg[63] ;
  reg \r_reg[32] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[32]  <= r_n[32];
  assign r[32] = \r_reg[32] ;
  reg \r_reg[33] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[33]  <= r_n[33];
  assign r[33] = \r_reg[33] ;
  reg \r_reg[34] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[34]  <= r_n[34];
  assign r[34] = \r_reg[34] ;
  reg \r_reg[35] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[35]  <= r_n[35];
  assign r[35] = \r_reg[35] ;
  reg \r_reg[36] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[36]  <= r_n[36];
  assign r[36] = \r_reg[36] ;
  reg \r_reg[37] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[37]  <= r_n[37];
  assign r[37] = \r_reg[37] ;
  reg \r_reg[38] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[38]  <= r_n[38];
  assign r[38] = \r_reg[38] ;
  reg \r_reg[39] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[39]  <= r_n[39];
  assign r[39] = \r_reg[39] ;
  reg \r_reg[40] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[40]  <= r_n[40];
  assign r[40] = \r_reg[40] ;
  reg \r_reg[41] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[41]  <= r_n[41];
  assign r[41] = \r_reg[41] ;
  reg \r_reg[42] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[42]  <= r_n[42];
  assign r[42] = \r_reg[42] ;
  reg \r_reg[43] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[43]  <= r_n[43];
  assign r[43] = \r_reg[43] ;
  reg \r_reg[44] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[44]  <= r_n[44];
  assign r[44] = \r_reg[44] ;
  reg \r_reg[45] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[45]  <= r_n[45];
  assign r[45] = \r_reg[45] ;
  reg \r_reg[46] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[46]  <= r_n[46];
  assign r[46] = \r_reg[46] ;
  reg \r_reg[47] ;
  always @(posedge clk_i)
    if (_0002_) \r_reg[47]  <= r_n[47];
  assign r[47] = \r_reg[47] ;
  reg \r_reg[16] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[16]  <= r_n[16];
  assign r[16] = \r_reg[16] ;
  reg \r_reg[17] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[17]  <= r_n[17];
  assign r[17] = \r_reg[17] ;
  reg \r_reg[18] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[18]  <= r_n[18];
  assign r[18] = \r_reg[18] ;
  reg \r_reg[19] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[19]  <= r_n[19];
  assign r[19] = \r_reg[19] ;
  reg \r_reg[20] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[20]  <= r_n[20];
  assign r[20] = \r_reg[20] ;
  reg \r_reg[21] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[21]  <= r_n[21];
  assign r[21] = \r_reg[21] ;
  reg \r_reg[22] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[22]  <= r_n[22];
  assign r[22] = \r_reg[22] ;
  reg \r_reg[23] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[23]  <= r_n[23];
  assign r[23] = \r_reg[23] ;
  reg \r_reg[24] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[24]  <= r_n[24];
  assign r[24] = \r_reg[24] ;
  reg \r_reg[25] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[25]  <= r_n[25];
  assign r[25] = \r_reg[25] ;
  reg \r_reg[26] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[26]  <= r_n[26];
  assign r[26] = \r_reg[26] ;
  reg \r_reg[27] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[27]  <= r_n[27];
  assign r[27] = \r_reg[27] ;
  reg \r_reg[28] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[28]  <= r_n[28];
  assign r[28] = \r_reg[28] ;
  reg \r_reg[29] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[29]  <= r_n[29];
  assign r[29] = \r_reg[29] ;
  reg \r_reg[30] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[30]  <= r_n[30];
  assign r[30] = \r_reg[30] ;
  reg \r_reg[31] ;
  always @(posedge clk_i)
    if (_0001_) \r_reg[31]  <= r_n[31];
  assign r[31] = \r_reg[31] ;
  reg \r_reg[496] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[496]  <= 1'h0;
      else \r_reg[496]  <= data_i[0];
  assign r[496] = \r_reg[496] ;
  reg \r_reg[497] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[497]  <= 1'h0;
      else \r_reg[497]  <= data_i[1];
  assign r[497] = \r_reg[497] ;
  reg \r_reg[498] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[498]  <= 1'h0;
      else \r_reg[498]  <= data_i[2];
  assign r[498] = \r_reg[498] ;
  reg \r_reg[499] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[499]  <= 1'h0;
      else \r_reg[499]  <= data_i[3];
  assign r[499] = \r_reg[499] ;
  reg \r_reg[500] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[500]  <= 1'h0;
      else \r_reg[500]  <= data_i[4];
  assign r[500] = \r_reg[500] ;
  reg \r_reg[501] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[501]  <= 1'h0;
      else \r_reg[501]  <= data_i[5];
  assign r[501] = \r_reg[501] ;
  reg \r_reg[502] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[502]  <= 1'h0;
      else \r_reg[502]  <= data_i[6];
  assign r[502] = \r_reg[502] ;
  reg \r_reg[503] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[503]  <= 1'h0;
      else \r_reg[503]  <= data_i[7];
  assign r[503] = \r_reg[503] ;
  reg \r_reg[504] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[504]  <= 1'h0;
      else \r_reg[504]  <= data_i[8];
  assign r[504] = \r_reg[504] ;
  reg \r_reg[505] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[505]  <= 1'h0;
      else \r_reg[505]  <= data_i[9];
  assign r[505] = \r_reg[505] ;
  reg \r_reg[506] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[506]  <= 1'h0;
      else \r_reg[506]  <= data_i[10];
  assign r[506] = \r_reg[506] ;
  reg \r_reg[507] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[507]  <= 1'h0;
      else \r_reg[507]  <= data_i[11];
  assign r[507] = \r_reg[507] ;
  reg \r_reg[508] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[508]  <= 1'h0;
      else \r_reg[508]  <= data_i[12];
  assign r[508] = \r_reg[508] ;
  reg \r_reg[509] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[509]  <= 1'h0;
      else \r_reg[509]  <= data_i[13];
  assign r[509] = \r_reg[509] ;
  reg \r_reg[510] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[510]  <= 1'h0;
      else \r_reg[510]  <= data_i[14];
  assign r[510] = \r_reg[510] ;
  reg \r_reg[511] ;
  always @(posedge clk_i)
    if (_0031_)
      if (_0032_) \r_reg[511]  <= 1'h0;
      else \r_reg[511]  <= data_i[15];
  assign r[511] = \r_reg[511] ;
  assign r[15:0] = data_o;
  assign r_n[511:496] = 16'hxxxx;
endmodule
