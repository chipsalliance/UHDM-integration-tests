module bsg_round_robin_n_to_1(clk_i, reset_i, data_i, v_i, yumi_o, v_o, data_o, tag_o, yumi_i);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  input clk_i;
  wire clk_i;
  input [31:0] data_i;
  wire [31:0] data_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire [1:0] \greedy.grants_lo ;
  wire \greedy.scan0.rr_arb_ctrl.clk_i ;
  wire \greedy.scan0.rr_arb_ctrl.grants_en_i ;
  wire [1:0] \greedy.scan0.rr_arb_ctrl.grants_o ;
  wire \greedy.scan0.rr_arb_ctrl.hold_on_sr ;
  wire [1:0] \greedy.scan0.rr_arb_ctrl.inputs_2.sel_one_hot_n ;
  reg \greedy.scan0.rr_arb_ctrl.last_r ;
  wire [1:0] \greedy.scan0.rr_arb_ctrl.reqs_i ;
  wire \greedy.scan0.rr_arb_ctrl.reset_i ;
  wire \greedy.scan0.rr_arb_ctrl.reset_on_sr ;
  wire [1:0] \greedy.scan0.rr_arb_ctrl.sel_one_hot_o ;
  wire \greedy.scan0.rr_arb_ctrl.tag_o ;
  wire \greedy.scan0.rr_arb_ctrl.v_o ;
  wire \greedy.scan0.rr_arb_ctrl.yumi_i ;
  wire [31:0] \greedy.xbar.i ;
  wire [31:0] \greedy.xbar.l[0].mux_one_hot.data_i ;
  wire [15:0] \greedy.xbar.l[0].mux_one_hot.data_o ;
  wire [1:0] \greedy.xbar.l[0].mux_one_hot.sel_one_hot_i ;
  wire [15:0] \greedy.xbar.o ;
  wire [1:0] \greedy.xbar.sel_oi_one_hot_i ;
  input reset_i;
  wire reset_i;
  output tag_o;
  wire tag_o;
  input [1:0] v_i;
  wire [1:0] v_i;
  output v_o;
  wire v_o;
  input yumi_i;
  wire yumi_i;
  output [1:0] yumi_o;
  wire [1:0] yumi_o;
  assign _013_ = ~v_i[0];
  assign _014_ = v_i[1] | ~(v_i[0]);
  assign _015_ = ~v_i[1];
  assign _016_ = v_i[0] | ~(v_i[1]);
  assign _017_ = \greedy.scan0.rr_arb_ctrl.last_r  ? _016_ : _015_;
  assign _018_ = \greedy.scan0.rr_arb_ctrl.last_r  ? _013_ : _014_;
  assign _019_ = data_i[0] & ~(_018_);
  assign _020_ = v_i[1] & ~(v_i[0]);
  assign \greedy.scan0.rr_arb_ctrl.tag_o  = \greedy.scan0.rr_arb_ctrl.last_r  ? _020_ : v_i[1];
  assign _021_ = _018_ & ~(\greedy.scan0.rr_arb_ctrl.tag_o );
  assign _022_ = _021_ | _017_;
  assign _023_ = data_i[16] & ~(_022_);
  assign data_o[0] = _023_ | _019_;
  assign _024_ = data_i[1] & ~(_018_);
  assign _025_ = data_i[17] & ~(_022_);
  assign data_o[1] = _025_ | _024_;
  assign _026_ = data_i[2] & ~(_018_);
  assign _027_ = data_i[18] & ~(_022_);
  assign data_o[2] = _027_ | _026_;
  assign _028_ = data_i[3] & ~(_018_);
  assign _029_ = data_i[19] & ~(_022_);
  assign data_o[3] = _029_ | _028_;
  assign _030_ = data_i[4] & ~(_018_);
  assign _031_ = data_i[20] & ~(_022_);
  assign data_o[4] = _031_ | _030_;
  assign _032_ = data_i[5] & ~(_018_);
  assign _033_ = data_i[21] & ~(_022_);
  assign data_o[5] = _033_ | _032_;
  assign _034_ = data_i[6] & ~(_018_);
  assign _035_ = data_i[22] & ~(_022_);
  assign data_o[6] = _035_ | _034_;
  assign _036_ = data_i[7] & ~(_018_);
  assign _037_ = data_i[23] & ~(_022_);
  assign data_o[7] = _037_ | _036_;
  assign _038_ = data_i[8] & ~(_018_);
  assign _039_ = data_i[24] & ~(_022_);
  assign data_o[8] = _039_ | _038_;
  assign _040_ = data_i[9] & ~(_018_);
  assign _041_ = data_i[25] & ~(_022_);
  assign data_o[9] = _041_ | _040_;
  assign _000_ = data_i[10] & ~(_018_);
  assign _001_ = data_i[26] & ~(_022_);
  assign data_o[10] = _001_ | _000_;
  assign _002_ = data_i[11] & ~(_018_);
  assign _003_ = data_i[27] & ~(_022_);
  assign data_o[11] = _003_ | _002_;
  assign _004_ = data_i[12] & ~(_018_);
  assign _005_ = data_i[28] & ~(_022_);
  assign data_o[12] = _005_ | _004_;
  assign _006_ = data_i[13] & ~(_018_);
  assign _007_ = data_i[29] & ~(_022_);
  assign data_o[13] = _007_ | _006_;
  assign _008_ = data_i[14] & ~(_018_);
  assign _009_ = data_i[30] & ~(_022_);
  assign data_o[14] = _009_ | _008_;
  assign _010_ = data_i[15] & ~(_018_);
  assign _011_ = data_i[31] & ~(_022_);
  assign data_o[15] = _011_ | _010_;
  assign _012_ = ~(v_i[1] | v_i[0]);
  assign v_o = ~_012_;
  assign yumi_o[0] = yumi_i & ~(_018_);
  assign yumi_o[1] = yumi_i & ~(_022_);
  assign \greedy.scan0.rr_arb_ctrl.yumi_i  = yumi_i & ~(_012_);
  always @(posedge clk_i)
    if (reset_i) \greedy.scan0.rr_arb_ctrl.last_r  <= 1'h0;
    else if (\greedy.scan0.rr_arb_ctrl.yumi_i ) \greedy.scan0.rr_arb_ctrl.last_r  <= \greedy.scan0.rr_arb_ctrl.tag_o ;
  assign \greedy.grants_lo  = \greedy.scan0.rr_arb_ctrl.grants_o ;
  assign \greedy.scan0.rr_arb_ctrl.clk_i  = clk_i;
  assign \greedy.scan0.rr_arb_ctrl.grants_en_i  = 1'h1;
  assign \greedy.scan0.rr_arb_ctrl.hold_on_sr  = 1'h0;
  assign \greedy.scan0.rr_arb_ctrl.inputs_2.sel_one_hot_n  = \greedy.scan0.rr_arb_ctrl.grants_o ;
  assign \greedy.scan0.rr_arb_ctrl.reqs_i  = v_i;
  assign \greedy.scan0.rr_arb_ctrl.reset_i  = reset_i;
  assign \greedy.scan0.rr_arb_ctrl.reset_on_sr  = 1'h0;
  assign \greedy.scan0.rr_arb_ctrl.sel_one_hot_o  = \greedy.scan0.rr_arb_ctrl.grants_o ;
  assign \greedy.scan0.rr_arb_ctrl.v_o  = v_o;
  assign \greedy.xbar.i  = data_i;
  assign \greedy.xbar.l[0].mux_one_hot.data_i  = data_i;
  assign \greedy.xbar.l[0].mux_one_hot.data_o  = data_o;
  assign \greedy.xbar.l[0].mux_one_hot.sel_one_hot_i  = \greedy.scan0.rr_arb_ctrl.grants_o ;
  assign \greedy.xbar.o  = data_o;
  assign \greedy.xbar.sel_oi_one_hot_i  = \greedy.scan0.rr_arb_ctrl.grants_o ;
  assign tag_o = \greedy.scan0.rr_arb_ctrl.tag_o ;
endmodule
