module bsg_dff_gatestack(i0, i1, o);
  input [15:0] i0;
  wire [15:0] i0;
  input [15:0] i1;
  wire [15:0] i1;
  output [15:0] o;
  reg [15:0] o;
  always @(posedge i1[15])
    o[15] <= i0[15];
  always @(posedge i1[14])
    o[14] <= i0[14];
  always @(posedge i1[13])
    o[13] <= i0[13];
  always @(posedge i1[12])
    o[12] <= i0[12];
  always @(posedge i1[11])
    o[11] <= i0[11];
  always @(posedge i1[10])
    o[10] <= i0[10];
  always @(posedge i1[9])
    o[9] <= i0[9];
  always @(posedge i1[8])
    o[8] <= i0[8];
  always @(posedge i1[7])
    o[7] <= i0[7];
  always @(posedge i1[6])
    o[6] <= i0[6];
  always @(posedge i1[5])
    o[5] <= i0[5];
  always @(posedge i1[4])
    o[4] <= i0[4];
  always @(posedge i1[3])
    o[3] <= i0[3];
  always @(posedge i1[2])
    o[2] <= i0[2];
  always @(posedge i1[1])
    o[1] <= i0[1];
  always @(posedge i1[0])
    o[0] <= i0[0];
endmodule
