module top;
  import flash_ctrl_pkg::*;
  logic [15:0] array [3];
  logic [2:0] q;
endmodule
