module bsg_round_robin_arb(clk_i, reset_i, grants_en_i, reqs_i, grants_o, sel_one_hot_o, v_o, tag_o, yumi_i);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  input clk_i;
  wire clk_i;
  input grants_en_i;
  wire grants_en_i;
  output [15:0] grants_o;
  wire [15:0] grants_o;
  wire hold_on_sr;
  wire [15:0] \inputs_16.sel_one_hot_n ;
  reg [3:0] last_r;
  input [15:0] reqs_i;
  wire [15:0] reqs_i;
  input reset_i;
  wire reset_i;
  wire reset_on_sr;
  output [15:0] sel_one_hot_o;
  wire [15:0] sel_one_hot_o;
  output [3:0] tag_o;
  wire [3:0] tag_o;
  output v_o;
  wire v_o;
  input yumi_i;
  wire yumi_i;
  assign _0747_ = reqs_i[1] | reqs_i[0];
  assign _0758_ = reqs_i[3] | reqs_i[2];
  assign _0769_ = _0758_ | _0747_;
  assign _0780_ = reqs_i[5] | reqs_i[4];
  assign _0791_ = reqs_i[7] | reqs_i[6];
  assign _0802_ = _0791_ | _0780_;
  assign _0813_ = _0802_ | _0769_;
  assign _0824_ = reqs_i[9] | reqs_i[8];
  assign _0835_ = reqs_i[11] | reqs_i[10];
  assign _0846_ = _0835_ | _0824_;
  assign _0857_ = reqs_i[13] | reqs_i[12];
  assign _0868_ = reqs_i[15] | reqs_i[14];
  assign _0879_ = _0868_ | _0857_;
  assign _0890_ = _0879_ | _0846_;
  assign v_o = _0890_ | _0813_;
  assign _0911_ = ~(reqs_i[0] & last_r[0]);
  assign _0922_ = ~(last_r[1] & last_r[2]);
  assign _0933_ = _0922_ | _0911_;
  assign _0944_ = last_r[3] & ~(_0933_);
  assign _0955_ = reqs_i[0] & ~(reqs_i[11]);
  assign _0966_ = _0955_ & ~(_0857_);
  assign _0977_ = last_r[0] | ~(last_r[1]);
  assign _0988_ = _0977_ | _0868_;
  assign _0999_ = _0966_ & ~(_0988_);
  assign _1010_ = last_r[2] | ~(last_r[3]);
  assign _1021_ = _0999_ & ~(_1010_);
  assign _1032_ = _1021_ | _0944_;
  assign _1043_ = reqs_i[0] & ~(reqs_i[10]);
  assign _1054_ = reqs_i[11] | reqs_i[12];
  assign _1065_ = _1043_ & ~(_1054_);
  assign _1076_ = reqs_i[13] | reqs_i[14];
  assign _1087_ = reqs_i[15] | ~(last_r[0]);
  assign _1098_ = _1087_ | _1076_;
  assign _1109_ = _1065_ & ~(_1098_);
  assign _1120_ = ~last_r[3];
  assign _1131_ = last_r[1] | last_r[2];
  assign _1142_ = _1131_ | _1120_;
  assign _1153_ = _1109_ & ~(_1142_);
  assign _1164_ = reqs_i[9] | ~(reqs_i[0]);
  assign _1175_ = _1164_ | _0835_;
  assign _1186_ = ~(_1175_ | _0879_);
  assign _0010_ = last_r[1] | last_r[0];
  assign _0021_ = _0010_ | _1010_;
  assign _0032_ = _1186_ & ~(_0021_);
  assign _0043_ = _0032_ | _1153_;
  assign _0054_ = _0043_ | _1032_;
  assign _0065_ = reqs_i[0] & ~(reqs_i[8]);
  assign _0076_ = reqs_i[9] | reqs_i[10];
  assign _0087_ = _0065_ & ~(_0076_);
  assign _0098_ = _1076_ | _1054_;
  assign _0109_ = _0087_ & ~(_0098_);
  assign _0120_ = _1087_ | _0922_;
  assign _0131_ = _0120_ | last_r[3];
  assign _0142_ = _0109_ & ~(_0131_);
  assign _0153_ = reqs_i[0] & ~(reqs_i[7]);
  assign _0164_ = _0153_ & ~(_0824_);
  assign _0175_ = _0857_ | _0835_;
  assign _0186_ = _0164_ & ~(_0175_);
  assign _0197_ = last_r[3] | ~(last_r[2]);
  assign _0208_ = _0197_ | _0988_;
  assign _0219_ = _0186_ & ~(_0208_);
  assign _0230_ = _0219_ | _0142_;
  assign _0241_ = reqs_i[0] & ~(reqs_i[6]);
  assign _0252_ = reqs_i[7] | reqs_i[8];
  assign _0256_ = _0241_ & ~(_0252_);
  assign _0258_ = _0076_ | _1054_;
  assign _0268_ = _0256_ & ~(_0258_);
  assign _0273_ = last_r[1] | ~(last_r[2]);
  assign _0274_ = _0273_ | last_r[3];
  assign _0275_ = _0274_ | _1098_;
  assign _0276_ = _0268_ & ~(_0275_);
  assign _0277_ = ~(_0835_ | _0824_);
  assign _0278_ = reqs_i[5] | ~(reqs_i[0]);
  assign _0279_ = _0278_ | _0791_;
  assign _0280_ = _0277_ & ~(_0279_);
  assign _0281_ = ~(last_r[1] | last_r[0]);
  assign _0282_ = _0281_ & ~(_0197_);
  assign _0283_ = _0879_ | ~(_0282_);
  assign _0284_ = _0280_ & ~(_0283_);
  assign _0285_ = _0284_ | _0276_;
  assign _0286_ = _0285_ | _0230_;
  assign _0287_ = _0286_ | _0054_;
  assign _0288_ = reqs_i[4] | ~(reqs_i[0]);
  assign _0289_ = reqs_i[5] | reqs_i[6];
  assign _0290_ = _0289_ | _0288_;
  assign _0291_ = _0252_ | _0076_;
  assign _0292_ = _0291_ | _0290_;
  assign _0293_ = last_r[2] | ~(last_r[1]);
  assign _0294_ = _0293_ | _1087_;
  assign _0295_ = _0294_ | _0098_;
  assign _0296_ = _0295_ | _0292_;
  assign _0297_ = _1120_ & ~(_0296_);
  assign _0298_ = reqs_i[0] & ~(reqs_i[3]);
  assign _0299_ = _0298_ & ~(_0780_);
  assign _0300_ = _0824_ | _0791_;
  assign _0301_ = _0299_ & ~(_0300_);
  assign _0302_ = _0175_ | _0988_;
  assign _0303_ = _0301_ & ~(_0302_);
  assign _0304_ = last_r[3] | last_r[2];
  assign _0305_ = _0303_ & ~(_0304_);
  assign _0306_ = _0305_ | _0297_;
  assign _0307_ = reqs_i[0] & ~(reqs_i[2]);
  assign _0308_ = reqs_i[3] | reqs_i[4];
  assign _0309_ = _0307_ & ~(_0308_);
  assign _0310_ = _0289_ | _0252_;
  assign _0311_ = _0309_ & ~(_0310_);
  assign _0312_ = _0258_ | _1098_;
  assign _0313_ = _0311_ & ~(_0312_);
  assign _0314_ = _1131_ | last_r[3];
  assign _0315_ = _0313_ & ~(_0314_);
  assign _0316_ = reqs_i[1] | ~(reqs_i[0]);
  assign _0317_ = _0316_ | _0758_;
  assign _0318_ = _0317_ | _0802_;
  assign _0319_ = ~(_0318_ | _0890_);
  assign _0320_ = _0304_ | _0010_;
  assign _0321_ = _0319_ & ~(_0320_);
  assign _0322_ = _0321_ | _0315_;
  assign _0323_ = _0322_ | _0306_;
  assign _0324_ = last_r[1] & ~(last_r[0]);
  assign _0325_ = reqs_i[15] | ~(reqs_i[0]);
  assign _0326_ = _0324_ & ~(_0325_);
  assign _0327_ = ~(last_r[3] & last_r[2]);
  assign _0328_ = _0326_ & ~(_0327_);
  assign _0329_ = reqs_i[0] & ~(reqs_i[14]);
  assign _0330_ = _0329_ & ~(_1087_);
  assign _0331_ = _0273_ | _1120_;
  assign _0332_ = _0330_ & ~(_0331_);
  assign _0333_ = _0332_ | _0328_;
  assign _0334_ = reqs_i[0] & ~(reqs_i[13]);
  assign _0335_ = _0334_ & ~(_0868_);
  assign _0336_ = _0327_ | _0010_;
  assign _0337_ = _0335_ & ~(_0336_);
  assign _0338_ = reqs_i[12] | ~(reqs_i[0]);
  assign _0339_ = _0338_ | _1076_;
  assign _0340_ = _0339_ | _0294_;
  assign _0341_ = last_r[3] & ~(_0340_);
  assign _0342_ = _0341_ | _0337_;
  assign _0343_ = _0342_ | _0333_;
  assign _0344_ = _0343_ | _0323_;
  assign _0345_ = _0344_ | _0287_;
  assign _0346_ = reqs_i[14] | ~(reqs_i[15]);
  assign _0347_ = _0346_ | _0857_;
  assign _0348_ = ~(_0347_ | _0846_);
  assign _0349_ = _0348_ & ~(_0813_);
  assign _0350_ = ~(last_r[1] & last_r[0]);
  assign _0351_ = _0350_ | _0327_;
  assign _0352_ = _0349_ & ~(_0351_);
  assign _0353_ = last_r[0] | ~(reqs_i[15]);
  assign _0354_ = _0353_ | _0293_;
  assign _0355_ = _0354_ | _0098_;
  assign _0356_ = last_r[3] & ~(_0355_);
  assign _0357_ = _0356_ | _0352_;
  assign _0358_ = last_r[3] & ~(last_r[2]);
  assign _0359_ = last_r[1] | ~(last_r[0]);
  assign _0360_ = _0359_ | _0346_;
  assign _0361_ = _0360_ | _0175_;
  assign _0362_ = _0358_ & ~(_0361_);
  assign _0363_ = ~_1142_;
  assign _0364_ = _0353_ | _1076_;
  assign _0365_ = _0364_ | _0258_;
  assign _0366_ = _0363_ & ~(_0365_);
  assign _0367_ = _0366_ | _0362_;
  assign _0368_ = _0367_ | _0357_;
  assign _0369_ = last_r[2] & ~(last_r[3]);
  assign _0370_ = _0350_ | ~(_0369_);
  assign _0371_ = _0348_ & ~(_0370_);
  assign _0372_ = ~(_1076_ | _1054_);
  assign _0373_ = _0372_ & ~(_0291_);
  assign _0374_ = _0353_ | _0922_;
  assign _0375_ = _0374_ | last_r[3];
  assign _0376_ = _0373_ & ~(_0375_);
  assign _0377_ = _0376_ | _0371_;
  assign _0378_ = ~(_0857_ | _0835_);
  assign _0379_ = _0378_ & ~(_0300_);
  assign _0380_ = _0360_ | ~(_0369_);
  assign _0381_ = _0379_ & ~(_0380_);
  assign _0382_ = ~(_0076_ | _1054_);
  assign _0383_ = _0382_ & ~(_0310_);
  assign _0384_ = _0364_ | _0274_;
  assign _0385_ = _0383_ & ~(_0384_);
  assign _0386_ = _0385_ | _0381_;
  assign _0387_ = _0386_ | _0377_;
  assign _0388_ = _0387_ | _0368_;
  assign _0389_ = _0277_ & ~(_0802_);
  assign _0390_ = ~(last_r[3] | last_r[2]);
  assign _0391_ = _0390_ & ~(_0350_);
  assign _0392_ = _0347_ | ~(_0391_);
  assign _0393_ = _0389_ & ~(_0392_);
  assign _0394_ = _0308_ | _0289_;
  assign _0395_ = ~(_0394_ | _0291_);
  assign _0396_ = _0355_ | ~(_0395_);
  assign _0397_ = _1120_ & ~(_0396_);
  assign _0398_ = _0397_ | _0393_;
  assign _0399_ = _0780_ | _0758_;
  assign _0400_ = _0399_ | _0300_;
  assign _0401_ = _0400_ | _0361_;
  assign _0402_ = _0390_ & ~(_0401_);
  assign _0403_ = ~_0314_;
  assign _0404_ = reqs_i[1] | reqs_i[2];
  assign _0405_ = _0404_ | _0308_;
  assign _0406_ = _0405_ | _0310_;
  assign _0407_ = _0406_ | _0365_;
  assign _0408_ = _0403_ & ~(_0407_);
  assign _0409_ = _0408_ | _0402_;
  assign _0410_ = _0409_ | _0398_;
  assign _0411_ = last_r[3] & ~(_0374_);
  assign _0412_ = ~(_0360_ | _0327_);
  assign _0413_ = _0412_ | _0411_;
  assign _0414_ = ~(_0364_ | _0331_);
  assign _0415_ = _0358_ & ~(_0350_);
  assign _0416_ = _0415_ & ~(_0347_);
  assign _0417_ = _0416_ | _0414_;
  assign _0418_ = _0417_ | _0413_;
  assign _0419_ = _0418_ | _0410_;
  assign _0420_ = _0419_ | _0388_;
  assign _0421_ = ~(last_r[0] & reqs_i[14]);
  assign _0422_ = _0421_ | _0857_;
  assign _0423_ = ~(_0422_ | _0846_);
  assign _0424_ = _0423_ & ~(_0813_);
  assign _0425_ = _0922_ | _1120_;
  assign _0426_ = _0424_ & ~(_0425_);
  assign _0427_ = ~(_0758_ | _0747_);
  assign _0428_ = _0427_ & ~(_0802_);
  assign _0429_ = reqs_i[15] | ~(reqs_i[14]);
  assign _0430_ = _0429_ | _0857_;
  assign _0431_ = _0430_ | _0846_;
  assign _0432_ = _0428_ & ~(_0431_);
  assign _0433_ = _0327_ | _0977_;
  assign _0434_ = _0432_ & ~(_0433_);
  assign _0435_ = _0434_ | _0426_;
  assign _0436_ = reqs_i[13] | ~(reqs_i[14]);
  assign _0437_ = _0436_ | _1054_;
  assign _0438_ = _0324_ & ~(_1010_);
  assign _0439_ = _0438_ & ~(_0437_);
  assign _0440_ = _0421_ | _1131_;
  assign _0441_ = _0440_ | _0175_;
  assign _0442_ = last_r[3] & ~(_0441_);
  assign _0443_ = _0442_ | _0439_;
  assign _0444_ = _0443_ | _0435_;
  assign _0445_ = _0436_ | _0010_;
  assign _0446_ = _0445_ | _0258_;
  assign _0447_ = _0358_ & ~(_0446_);
  assign _0448_ = _0922_ | last_r[3];
  assign _0449_ = _0423_ & ~(_0448_);
  assign _0450_ = _0449_ | _0447_;
  assign _0451_ = ~(_0437_ | _0291_);
  assign _0452_ = _0197_ | _0977_;
  assign _0453_ = _0451_ & ~(_0452_);
  assign _0454_ = _0421_ | _0273_;
  assign _0455_ = _0454_ | last_r[3];
  assign _0456_ = _0379_ & ~(_0455_);
  assign _0457_ = _0456_ | _0453_;
  assign _0458_ = _0457_ | _0450_;
  assign _0459_ = _0458_ | _0444_;
  assign _0460_ = _0445_ | ~(_0369_);
  assign _0461_ = _0383_ & ~(_0460_);
  assign _0462_ = _0293_ | last_r[3];
  assign _0463_ = _0462_ | _0422_;
  assign _0464_ = _0389_ & ~(_0463_);
  assign _0465_ = _0464_ | _0461_;
  assign _0466_ = _0324_ & ~(_0304_);
  assign _0467_ = _0437_ | ~(_0466_);
  assign _0468_ = _0395_ & ~(_0467_);
  assign _0469_ = _0441_ | _0400_;
  assign _0470_ = _1120_ & ~(_0469_);
  assign _0471_ = _0470_ | _0468_;
  assign _0472_ = _0471_ | _0465_;
  assign _0473_ = _0446_ | _0406_;
  assign _0474_ = _0390_ & ~(_0473_);
  assign _0475_ = last_r[3] & ~(_0454_);
  assign _0476_ = _0475_ | _0474_;
  assign _0477_ = ~(_0445_ | _0327_);
  assign _0478_ = _0293_ | _1120_;
  assign _0479_ = ~(_0478_ | _0422_);
  assign _0480_ = _0479_ | _0477_;
  assign _0481_ = _0480_ | _0476_;
  assign _0482_ = _0481_ | _0472_;
  assign _0483_ = _0482_ | _0459_;
  assign _0484_ = ~(_0483_ | _0420_);
  assign _0485_ = reqs_i[12] | ~(reqs_i[13]);
  assign _0486_ = _0485_ | _0350_;
  assign _0487_ = _0486_ | _0846_;
  assign _0488_ = _0487_ | _0813_;
  assign _0489_ = ~(_0488_ | _0327_);
  assign _0490_ = ~_0425_;
  assign _0491_ = last_r[0] | reqs_i[15];
  assign _0492_ = _0491_ | _0485_;
  assign _0493_ = _0492_ | _0846_;
  assign _0494_ = _0493_ | _0813_;
  assign _0495_ = _0490_ & ~(_0494_);
  assign _0496_ = _0495_ | _0489_;
  assign _0497_ = last_r[0] | ~(reqs_i[13]);
  assign _0498_ = _0497_ | _1054_;
  assign _0499_ = ~(_0498_ | _0478_);
  assign _0500_ = _0485_ | _0835_;
  assign _0501_ = _0358_ & ~(_0359_);
  assign _0502_ = _0501_ & ~(_0500_);
  assign _0503_ = _0502_ | _0499_;
  assign _0504_ = _0503_ | _0496_;
  assign _0505_ = _0497_ | _1131_;
  assign _0506_ = _0505_ | _0258_;
  assign _0507_ = last_r[3] & ~(_0506_);
  assign _0508_ = _0369_ & ~(_0487_);
  assign _0509_ = _0508_ | _0507_;
  assign _0510_ = ~_0448_;
  assign _0511_ = _0498_ | _0291_;
  assign _0512_ = _0510_ & ~(_0511_);
  assign _0513_ = ~(_0500_ | _0300_);
  assign _0514_ = _0359_ | ~(_0369_);
  assign _0515_ = _0513_ & ~(_0514_);
  assign _0516_ = _0515_ | _0512_;
  assign _0517_ = _0516_ | _0509_;
  assign _0518_ = _0517_ | _0504_;
  assign _0519_ = _0497_ | _0273_;
  assign _0520_ = _0519_ | last_r[3];
  assign _0521_ = _0383_ & ~(_0520_);
  assign _0522_ = _0486_ | ~(_0390_);
  assign _0523_ = _0389_ & ~(_0522_);
  assign _0524_ = _0523_ | _0521_;
  assign _0525_ = _0498_ | _0462_;
  assign _0526_ = _0395_ & ~(_0525_);
  assign _0527_ = ~(_0399_ | _0300_);
  assign _0528_ = _0390_ & ~(_0359_);
  assign _0529_ = _0500_ | ~(_0528_);
  assign _0530_ = _0527_ & ~(_0529_);
  assign _0531_ = _0530_ | _0526_;
  assign _0532_ = _0531_ | _0524_;
  assign _0533_ = _0506_ | _0406_;
  assign _0534_ = _1120_ & ~(_0533_);
  assign _0535_ = _0485_ | _0868_;
  assign _0536_ = _0535_ | _0846_;
  assign _0537_ = ~(_0536_ | _0813_);
  assign _0538_ = _0359_ | _0327_;
  assign _0539_ = _0537_ & ~(_0538_);
  assign _0540_ = _0539_ | _0534_;
  assign _0541_ = last_r[3] & ~(_0519_);
  assign _0542_ = _0358_ & ~(_0486_);
  assign _0543_ = _0542_ | _0541_;
  assign _0544_ = _0543_ | _0540_;
  assign _0545_ = _0544_ | _0532_;
  assign _0546_ = _0545_ | _0518_;
  assign _0547_ = ~(last_r[0] & reqs_i[12]);
  assign _0548_ = _0547_ | _0922_;
  assign _0549_ = _0548_ | _0846_;
  assign _0550_ = _0549_ | _0813_;
  assign _0551_ = last_r[3] & ~(_0550_);
  assign _0552_ = reqs_i[11] | ~(reqs_i[12]);
  assign _0553_ = _0552_ | _0977_;
  assign _0554_ = _0358_ & ~(_0553_);
  assign _0555_ = _0554_ | _0551_;
  assign _0556_ = _0547_ | _0835_;
  assign _0557_ = ~(_0556_ | _1142_);
  assign _0558_ = _0552_ | _0076_;
  assign _0559_ = ~(_0558_ | _0021_);
  assign _0560_ = _0559_ | _0557_;
  assign _0561_ = _0560_ | _0555_;
  assign _0562_ = _1120_ & ~(_0549_);
  assign _0563_ = _0553_ | _0291_;
  assign _0564_ = _0369_ & ~(_0563_);
  assign _0565_ = _0564_ | _0562_;
  assign _0566_ = ~_0274_;
  assign _0567_ = _0556_ | _0300_;
  assign _0568_ = _0566_ & ~(_0567_);
  assign _0569_ = _0558_ | _0310_;
  assign _0570_ = _0282_ & ~(_0569_);
  assign _0571_ = _0570_ | _0568_;
  assign _0572_ = _0571_ | _0565_;
  assign _0573_ = _0572_ | _0561_;
  assign _0574_ = _0547_ | _0293_;
  assign _0575_ = _0574_ | last_r[3];
  assign _0576_ = _0389_ & ~(_0575_);
  assign _0577_ = _0553_ | _0304_;
  assign _0578_ = _0395_ & ~(_0577_);
  assign _0579_ = _0578_ | _0576_;
  assign _0580_ = _0556_ | _0314_;
  assign _0581_ = _0527_ & ~(_0580_);
  assign _0582_ = ~(_0405_ | _0310_);
  assign _0583_ = _0558_ | _0320_;
  assign _0584_ = _0582_ & ~(_0583_);
  assign _0585_ = _0584_ | _0581_;
  assign _0586_ = _0585_ | _0579_;
  assign _0587_ = ~_0327_;
  assign _0588_ = reqs_i[15] | ~(reqs_i[12]);
  assign _0589_ = _0588_ | _0977_;
  assign _0590_ = _0589_ | _0846_;
  assign _0591_ = _0590_ | _0813_;
  assign _0592_ = _0587_ & ~(_0591_);
  assign _0593_ = ~_0331_;
  assign _0594_ = reqs_i[14] | ~(reqs_i[12]);
  assign _0595_ = _0594_ | _1087_;
  assign _0596_ = _0595_ | _0846_;
  assign _0597_ = _0596_ | _0813_;
  assign _0598_ = _0593_ & ~(_0597_);
  assign _0599_ = _0598_ | _0592_;
  assign _0600_ = ~_0336_;
  assign _0601_ = reqs_i[13] | ~(reqs_i[12]);
  assign _0602_ = _0601_ | _0868_;
  assign _0603_ = _0602_ | _0846_;
  assign _0604_ = _0603_ | _0813_;
  assign _0605_ = _0600_ & ~(_0604_);
  assign _0606_ = last_r[3] & ~(_0574_);
  assign _0607_ = _0606_ | _0605_;
  assign _0608_ = _0607_ | _0599_;
  assign _0609_ = _0608_ | _0586_;
  assign _0610_ = _0609_ | _0573_;
  assign _0611_ = _0610_ | _0546_;
  assign _0612_ = _0484_ & ~(_0611_);
  assign _0613_ = reqs_i[10] | ~(reqs_i[11]);
  assign _0614_ = _0613_ | _0824_;
  assign _0615_ = _0614_ | _0351_;
  assign _0616_ = ~(_0615_ | _0813_);
  assign _0617_ = last_r[0] | ~(reqs_i[11]);
  assign _0618_ = _0617_ | _0293_;
  assign _0619_ = last_r[3] & ~(_0618_);
  assign _0620_ = _0619_ | _0616_;
  assign _0621_ = _0613_ | _0359_;
  assign _0622_ = _0358_ & ~(_0621_);
  assign _0623_ = _0617_ | _0076_;
  assign _0624_ = ~(_0623_ | _1142_);
  assign _0625_ = _0624_ | _0622_;
  assign _0626_ = _0625_ | _0620_;
  assign _0627_ = ~(_0614_ | _0370_);
  assign _0628_ = _0617_ | _0922_;
  assign _0629_ = _0628_ | _0291_;
  assign _0630_ = _1120_ & ~(_0629_);
  assign _0631_ = _0630_ | _0627_;
  assign _0632_ = _0621_ | _0300_;
  assign _0633_ = _0369_ & ~(_0632_);
  assign _0634_ = _0623_ | _0310_;
  assign _0635_ = _0566_ & ~(_0634_);
  assign _0636_ = _0635_ | _0633_;
  assign _0637_ = _0636_ | _0631_;
  assign _0638_ = _0637_ | _0626_;
  assign _0639_ = _0614_ | _0802_;
  assign _0640_ = _0391_ & ~(_0639_);
  assign _0641_ = _0618_ | last_r[3];
  assign _0642_ = _0395_ & ~(_0641_);
  assign _0643_ = _0642_ | _0640_;
  assign _0644_ = _0621_ | _0304_;
  assign _0645_ = _0527_ & ~(_0644_);
  assign _0646_ = _0623_ | _0314_;
  assign _0647_ = _0582_ & ~(_0646_);
  assign _0648_ = _0647_ | _0645_;
  assign _0649_ = _0648_ | _0643_;
  assign _0650_ = _0491_ | _0922_;
  assign _0651_ = _0650_ | _0614_;
  assign _0652_ = _0651_ | _0813_;
  assign _0653_ = last_r[3] & ~(_0652_);
  assign _0654_ = _0359_ | _0868_;
  assign _0655_ = _0654_ | _0614_;
  assign _0656_ = _0655_ | _0813_;
  assign _0657_ = _0587_ & ~(_0656_);
  assign _0658_ = _0657_ | _0653_;
  assign _0659_ = _0491_ | _1076_;
  assign _0660_ = _0659_ | _0614_;
  assign _0661_ = _0660_ | _0813_;
  assign _0662_ = _0593_ & ~(_0661_);
  assign _0663_ = _0614_ | _0879_;
  assign _0664_ = _0663_ | _0813_;
  assign _0665_ = _0415_ & ~(_0664_);
  assign _0666_ = _0665_ | _0662_;
  assign _0667_ = _0666_ | _0658_;
  assign _0668_ = _0667_ | _0649_;
  assign _0669_ = _0668_ | _0638_;
  assign _0670_ = ~(last_r[0] & reqs_i[10]);
  assign _0671_ = _0670_ | _0824_;
  assign _0672_ = _0671_ | _0425_;
  assign _0673_ = ~(_0672_ | _0813_);
  assign _0674_ = _0670_ | _1131_;
  assign _0675_ = last_r[3] & ~(_0674_);
  assign _0676_ = _0675_ | _0673_;
  assign _0677_ = reqs_i[9] | ~(reqs_i[10]);
  assign _0678_ = _0677_ | _0010_;
  assign _0679_ = _0358_ & ~(_0678_);
  assign _0680_ = ~(_0671_ | _0448_);
  assign _0681_ = _0680_ | _0679_;
  assign _0682_ = _0681_ | _0676_;
  assign _0683_ = _0677_ | _0252_;
  assign _0684_ = ~(_0683_ | _0452_);
  assign _0685_ = _0670_ | _0273_;
  assign _0686_ = _0685_ | _0300_;
  assign _0687_ = _1120_ & ~(_0686_);
  assign _0688_ = _0687_ | _0684_;
  assign _0689_ = _0678_ | _0310_;
  assign _0690_ = _0369_ & ~(_0689_);
  assign _0691_ = ~_0462_;
  assign _0692_ = _0671_ | _0802_;
  assign _0693_ = _0691_ & ~(_0692_);
  assign _0694_ = _0693_ | _0690_;
  assign _0695_ = _0694_ | _0688_;
  assign _0696_ = _0695_ | _0682_;
  assign _0697_ = _0683_ | _0394_;
  assign _0698_ = _0466_ & ~(_0697_);
  assign _0699_ = _0674_ | last_r[3];
  assign _0700_ = _0527_ & ~(_0699_);
  assign _0701_ = _0700_ | _0698_;
  assign _0702_ = _0678_ | _0304_;
  assign _0703_ = _0582_ & ~(_0702_);
  assign _0704_ = reqs_i[15] | ~(reqs_i[10]);
  assign _0705_ = _0704_ | _0824_;
  assign _0706_ = _0705_ | _0433_;
  assign _0707_ = _0428_ & ~(_0706_);
  assign _0708_ = _0707_ | _0703_;
  assign _0709_ = _0708_ | _0701_;
  assign _0710_ = reqs_i[14] | ~(reqs_i[10]);
  assign _0711_ = _0710_ | _0824_;
  assign _0712_ = _0273_ | _1087_;
  assign _0713_ = _0712_ | _0711_;
  assign _0714_ = _0713_ | _0813_;
  assign _0715_ = last_r[3] & ~(_0714_);
  assign _0716_ = reqs_i[13] | ~(reqs_i[10]);
  assign _0717_ = _0716_ | _0824_;
  assign _0718_ = _0010_ | _0868_;
  assign _0719_ = _0718_ | _0717_;
  assign _0720_ = _0719_ | _0813_;
  assign _0721_ = _0587_ & ~(_0720_);
  assign _0722_ = _0721_ | _0715_;
  assign _0723_ = ~_0478_;
  assign _0724_ = reqs_i[12] | ~(reqs_i[10]);
  assign _0725_ = _0724_ | _0824_;
  assign _0726_ = _0725_ | _1098_;
  assign _0727_ = _0726_ | _0813_;
  assign _0728_ = _0723_ & ~(_0727_);
  assign _0729_ = reqs_i[11] | ~(reqs_i[10]);
  assign _0730_ = _0729_ | _0824_;
  assign _0731_ = _0730_ | _0879_;
  assign _0732_ = _0731_ | _0813_;
  assign _0733_ = _0438_ & ~(_0732_);
  assign _0734_ = _0733_ | _0728_;
  assign _0735_ = _0734_ | _0722_;
  assign _0736_ = _0735_ | _0709_;
  assign _0737_ = _0736_ | _0696_;
  assign _0738_ = _0737_ | _0669_;
  assign _0739_ = reqs_i[8] | ~(reqs_i[9]);
  assign _0740_ = _0739_ | _0350_;
  assign _0741_ = _0740_ | _0327_;
  assign _0742_ = ~(_0741_ | _0813_);
  assign _0743_ = _0739_ | _0835_;
  assign _0744_ = _0743_ | _0879_;
  assign _0745_ = _0744_ | _0813_;
  assign _0746_ = _0501_ & ~(_0745_);
  assign _0748_ = _0746_ | _0742_;
  assign _0749_ = last_r[0] | ~(reqs_i[9]);
  assign _0750_ = _0749_ | _1131_;
  assign _0751_ = last_r[3] & ~(_0750_);
  assign _0752_ = _0369_ & ~(_0740_);
  assign _0753_ = _0752_ | _0751_;
  assign _0754_ = _0753_ | _0748_;
  assign _0755_ = _0749_ | _0252_;
  assign _0756_ = ~(_0755_ | _0448_);
  assign _0757_ = _0739_ | _0791_;
  assign _0759_ = ~(_0757_ | _0514_);
  assign _0760_ = _0759_ | _0756_;
  assign _0761_ = _0749_ | _0273_;
  assign _0762_ = _0761_ | _0310_;
  assign _0763_ = _1120_ & ~(_0762_);
  assign _0764_ = _0740_ | _0802_;
  assign _0765_ = _0390_ & ~(_0764_);
  assign _0766_ = _0765_ | _0763_;
  assign _0767_ = _0766_ | _0760_;
  assign _0768_ = _0767_ | _0754_;
  assign _0770_ = _0755_ | _0394_;
  assign _0771_ = _0691_ & ~(_0770_);
  assign _0772_ = _0757_ | _0399_;
  assign _0773_ = _0528_ & ~(_0772_);
  assign _0774_ = _0773_ | _0771_;
  assign _0775_ = _0750_ | last_r[3];
  assign _0776_ = _0582_ & ~(_0775_);
  assign _0777_ = _0739_ | _0491_;
  assign _0778_ = _0777_ | _0425_;
  assign _0779_ = _0428_ & ~(_0778_);
  assign _0781_ = _0779_ | _0776_;
  assign _0782_ = _0781_ | _0774_;
  assign _0783_ = _0739_ | _0868_;
  assign _0784_ = _0783_ | _0538_;
  assign _0785_ = _0428_ & ~(_0784_);
  assign _0786_ = _0739_ | _1076_;
  assign _0787_ = _0491_ | _0273_;
  assign _0788_ = _0787_ | _0786_;
  assign _0789_ = _0788_ | _0813_;
  assign _0790_ = last_r[3] & ~(_0789_);
  assign _0792_ = _0790_ | _0785_;
  assign _0793_ = _0739_ | _0857_;
  assign _0794_ = _0350_ | _0868_;
  assign _0795_ = _0794_ | _0793_;
  assign _0796_ = _0795_ | _0813_;
  assign _0797_ = _0358_ & ~(_0796_);
  assign _0798_ = _0739_ | _1054_;
  assign _0799_ = _0798_ | _0659_;
  assign _0800_ = _0799_ | _0813_;
  assign _0801_ = _0723_ & ~(_0800_);
  assign _0803_ = _0801_ | _0797_;
  assign _0804_ = _0803_ | _0792_;
  assign _0805_ = _0804_ | _0782_;
  assign _0806_ = _0805_ | _0768_;
  assign _0807_ = ~(reqs_i[8] & last_r[0]);
  assign _0808_ = _0807_ | _0922_;
  assign _0809_ = _0808_ | _1120_;
  assign _0810_ = ~(_0809_ | _0813_);
  assign _0811_ = reqs_i[10] | ~(reqs_i[8]);
  assign _0812_ = _0811_ | _1054_;
  assign _0814_ = _0812_ | _1098_;
  assign _0815_ = _0814_ | _0813_;
  assign _0816_ = _0363_ & ~(_0815_);
  assign _0817_ = _0816_ | _0810_;
  assign _0818_ = reqs_i[9] | ~(reqs_i[8]);
  assign _0819_ = _0818_ | _0835_;
  assign _0820_ = _0819_ | _0879_;
  assign _0821_ = ~(_0820_ | _0813_);
  assign _0822_ = _0821_ & ~(_0021_);
  assign _0823_ = _1120_ & ~(_0808_);
  assign _0825_ = _0823_ | _0822_;
  assign _0826_ = _0825_ | _0817_;
  assign _0827_ = reqs_i[7] | ~(reqs_i[8]);
  assign _0828_ = _0827_ | _0977_;
  assign _0829_ = _0369_ & ~(_0828_);
  assign _0830_ = _0807_ | _0791_;
  assign _0831_ = ~(_0830_ | _0274_);
  assign _0832_ = _0831_ | _0829_;
  assign _0833_ = _0827_ | _0289_;
  assign _0834_ = _0282_ & ~(_0833_);
  assign _0836_ = _0807_ | _0293_;
  assign _0837_ = _0836_ | _0802_;
  assign _0838_ = _1120_ & ~(_0837_);
  assign _0839_ = _0838_ | _0834_;
  assign _0840_ = _0839_ | _0832_;
  assign _0841_ = _0840_ | _0826_;
  assign _0842_ = _0828_ | _0394_;
  assign _0843_ = _0390_ & ~(_0842_);
  assign _0844_ = _0830_ | _0399_;
  assign _0845_ = _0403_ & ~(_0844_);
  assign _0847_ = _0845_ | _0843_;
  assign _0848_ = ~_0320_;
  assign _0849_ = _0833_ | _0405_;
  assign _0850_ = _0848_ & ~(_0849_);
  assign _0851_ = reqs_i[15] | ~(reqs_i[8]);
  assign _0852_ = _0851_ | _0977_;
  assign _0853_ = _0852_ | _0327_;
  assign _0854_ = _0428_ & ~(_0853_);
  assign _0855_ = _0854_ | _0850_;
  assign _0856_ = _0855_ | _0847_;
  assign _0858_ = reqs_i[14] | ~(reqs_i[8]);
  assign _0859_ = _0858_ | _1087_;
  assign _0860_ = _0859_ | _0331_;
  assign _0861_ = _0428_ & ~(_0860_);
  assign _0862_ = reqs_i[13] | ~(reqs_i[8]);
  assign _0863_ = _0862_ | _0868_;
  assign _0864_ = _0863_ | _0336_;
  assign _0865_ = _0428_ & ~(_0864_);
  assign _0866_ = _0865_ | _0861_;
  assign _0867_ = reqs_i[12] | ~(reqs_i[8]);
  assign _0869_ = _0867_ | _1076_;
  assign _0870_ = _0869_ | _0294_;
  assign _0871_ = _0870_ | _0813_;
  assign _0872_ = last_r[3] & ~(_0871_);
  assign _0873_ = reqs_i[11] | ~(reqs_i[8]);
  assign _0874_ = _0873_ | _0857_;
  assign _0875_ = _0874_ | _0988_;
  assign _0876_ = _0875_ | _0813_;
  assign _0877_ = _0358_ & ~(_0876_);
  assign _0878_ = _0877_ | _0872_;
  assign _0880_ = _0878_ | _0866_;
  assign _0881_ = _0880_ | _0856_;
  assign _0882_ = _0881_ | _0841_;
  assign _0883_ = _0882_ | _0806_;
  assign _0884_ = _0883_ | _0738_;
  assign _0885_ = _0612_ & ~(_0884_);
  assign _0886_ = reqs_i[6] | ~(reqs_i[7]);
  assign _0887_ = _0886_ | _0780_;
  assign _0888_ = _0887_ | _0769_;
  assign _0889_ = ~(_0888_ | _0351_);
  assign _0891_ = _0654_ | _0175_;
  assign _0892_ = _0891_ | _0888_;
  assign _0893_ = _0358_ & ~(_0892_);
  assign _0894_ = _0893_ | _0889_;
  assign _0895_ = _0659_ | _0258_;
  assign _0896_ = _0895_ | _0888_;
  assign _0897_ = _0363_ & ~(_0896_);
  assign _0898_ = ~(_0887_ | _0769_);
  assign _0899_ = _0898_ & ~(_0890_);
  assign _0900_ = _0899_ & ~(_0370_);
  assign _0901_ = _0900_ | _0897_;
  assign _0902_ = _0901_ | _0894_;
  assign _0903_ = last_r[0] | ~(reqs_i[7]);
  assign _0904_ = _0903_ | _0922_;
  assign _0905_ = _1120_ & ~(_0904_);
  assign _0906_ = _0886_ | _0359_;
  assign _0907_ = _0369_ & ~(_0906_);
  assign _0908_ = _0907_ | _0905_;
  assign _0909_ = _0903_ | _0289_;
  assign _0910_ = ~(_0909_ | _0274_);
  assign _0912_ = _0391_ & ~(_0887_);
  assign _0913_ = _0912_ | _0910_;
  assign _0914_ = _0913_ | _0908_;
  assign _0915_ = _0914_ | _0902_;
  assign _0916_ = _0903_ | _0293_;
  assign _0917_ = _0916_ | _0394_;
  assign _0918_ = _1120_ & ~(_0917_);
  assign _0919_ = _0906_ | _0399_;
  assign _0920_ = _0390_ & ~(_0919_);
  assign _0921_ = _0920_ | _0918_;
  assign _0923_ = _0909_ | _0405_;
  assign _0924_ = _0403_ & ~(_0923_);
  assign _0925_ = _0650_ | _1120_;
  assign _0926_ = _0898_ & ~(_0925_);
  assign _0927_ = _0926_ | _0924_;
  assign _0928_ = _0927_ | _0921_;
  assign _0929_ = _0654_ | _0327_;
  assign _0930_ = _0898_ & ~(_0929_);
  assign _0931_ = _0659_ | _0331_;
  assign _0932_ = _0898_ & ~(_0931_);
  assign _0934_ = _0932_ | _0930_;
  assign _0935_ = _0879_ | ~(_0415_);
  assign _0936_ = _0898_ & ~(_0935_);
  assign _0937_ = _0491_ | _0293_;
  assign _0938_ = _0937_ | _0098_;
  assign _0939_ = _0938_ | _0888_;
  assign _0940_ = last_r[3] & ~(_0939_);
  assign _0941_ = _0940_ | _0936_;
  assign _0942_ = _0941_ | _0934_;
  assign _0943_ = _0942_ | _0928_;
  assign _0945_ = _0943_ | _0915_;
  assign _0946_ = ~(reqs_i[6] & last_r[0]);
  assign _0947_ = _0946_ | _0780_;
  assign _0948_ = _0947_ | _0769_;
  assign _0949_ = ~(_0948_ | _0425_);
  assign _0950_ = reqs_i[10] | ~(reqs_i[6]);
  assign _0951_ = _0950_ | _0780_;
  assign _0952_ = _0951_ | _0769_;
  assign _0953_ = _1131_ | _1087_;
  assign _0954_ = _0953_ | _0098_;
  assign _0956_ = _0954_ | _0952_;
  assign _0957_ = last_r[3] & ~(_0956_);
  assign _0958_ = _0957_ | _0949_;
  assign _0959_ = reqs_i[9] | ~(reqs_i[6]);
  assign _0960_ = _0959_ | _0780_;
  assign _0961_ = _0960_ | _0769_;
  assign _0962_ = _0718_ | _0175_;
  assign _0963_ = _0962_ | _0961_;
  assign _0964_ = _0358_ & ~(_0963_);
  assign _0965_ = reqs_i[8] | ~(reqs_i[6]);
  assign _0967_ = _0965_ | _0780_;
  assign _0968_ = _0967_ | _0769_;
  assign _0969_ = _0968_ | _0312_;
  assign _0970_ = _0510_ & ~(_0969_);
  assign _0971_ = _0970_ | _0964_;
  assign _0972_ = _0971_ | _0958_;
  assign _0973_ = reqs_i[7] | ~(reqs_i[6]);
  assign _0974_ = _0973_ | _0780_;
  assign _0975_ = _0974_ | _0769_;
  assign _0976_ = ~(_0975_ | _0890_);
  assign _0978_ = _0976_ & ~(_0452_);
  assign _0979_ = _0946_ | _0273_;
  assign _0980_ = _1120_ & ~(_0979_);
  assign _0981_ = _0980_ | _0978_;
  assign _0982_ = reqs_i[5] | ~(reqs_i[6]);
  assign _0983_ = _0982_ | _0010_;
  assign _0984_ = _0369_ & ~(_0983_);
  assign _0985_ = ~(_0947_ | _0462_);
  assign _0986_ = _0985_ | _0984_;
  assign _0987_ = _0986_ | _0981_;
  assign _0989_ = _0987_ | _0972_;
  assign _0990_ = _0982_ | _0308_;
  assign _0991_ = _0466_ & ~(_0990_);
  assign _0992_ = _0946_ | _1131_;
  assign _0993_ = _0992_ | _0399_;
  assign _0994_ = _1120_ & ~(_0993_);
  assign _0995_ = _0994_ | _0991_;
  assign _0996_ = _0983_ | _0405_;
  assign _0997_ = _0390_ & ~(_0996_);
  assign _0998_ = ~_0433_;
  assign _1000_ = reqs_i[15] | ~(reqs_i[6]);
  assign _1001_ = _1000_ | _0780_;
  assign _1002_ = _1001_ | _0769_;
  assign _1003_ = _0998_ & ~(_1002_);
  assign _1004_ = _1003_ | _0997_;
  assign _1005_ = _1004_ | _0995_;
  assign _1006_ = reqs_i[14] | ~(reqs_i[6]);
  assign _1007_ = _1006_ | _0780_;
  assign _1008_ = _0427_ & ~(_1007_);
  assign _1009_ = _0712_ | _1120_;
  assign _1011_ = _1008_ & ~(_1009_);
  assign _1012_ = reqs_i[13] | ~(reqs_i[6]);
  assign _1013_ = _1012_ | _0780_;
  assign _1014_ = _0427_ & ~(_1013_);
  assign _1015_ = _0718_ | _0327_;
  assign _1016_ = _1014_ & ~(_1015_);
  assign _1017_ = _1016_ | _1011_;
  assign _1018_ = reqs_i[12] | ~(reqs_i[6]);
  assign _1019_ = _1018_ | _0780_;
  assign _1020_ = _0427_ & ~(_1019_);
  assign _1022_ = _0478_ | _1098_;
  assign _1023_ = _1020_ & ~(_1022_);
  assign _1024_ = reqs_i[11] | ~(reqs_i[6]);
  assign _1025_ = _1024_ | _0780_;
  assign _1026_ = _0427_ & ~(_1025_);
  assign _1027_ = _0879_ | ~(_0438_);
  assign _1028_ = _1026_ & ~(_1027_);
  assign _1029_ = _1028_ | _1023_;
  assign _1030_ = _1029_ | _1017_;
  assign _1031_ = _1030_ | _1005_;
  assign _1033_ = _1031_ | _0989_;
  assign _1034_ = _1033_ | _0945_;
  assign _1035_ = reqs_i[4] | ~(reqs_i[5]);
  assign _1036_ = _1035_ | _0350_;
  assign _1037_ = _1036_ | _0769_;
  assign _1038_ = ~(_1037_ | _0327_);
  assign _1039_ = _1035_ | _0835_;
  assign _1040_ = _0427_ & ~(_1039_);
  assign _1041_ = _0879_ | ~(_0501_);
  assign _1042_ = _1040_ & ~(_1041_);
  assign _1044_ = _1042_ | _1038_;
  assign _1045_ = _1035_ | _0076_;
  assign _1046_ = _1045_ | _0769_;
  assign _1047_ = _0491_ | _1131_;
  assign _1048_ = _1047_ | _0098_;
  assign _1049_ = _1048_ | _1046_;
  assign _1050_ = last_r[3] & ~(_1049_);
  assign _1051_ = _1035_ | _0824_;
  assign _1052_ = _1051_ | _0769_;
  assign _1053_ = _0794_ | _0175_;
  assign _1055_ = _1053_ | _1052_;
  assign _1056_ = _0369_ & ~(_1055_);
  assign _1057_ = _1056_ | _1050_;
  assign _1058_ = _1057_ | _1044_;
  assign _1059_ = _1035_ | _0252_;
  assign _1060_ = _1059_ | _0769_;
  assign _1061_ = _1060_ | _0895_;
  assign _1062_ = _0510_ & ~(_1061_);
  assign _1063_ = _1035_ | _0791_;
  assign _1064_ = _1063_ | _0769_;
  assign _1066_ = ~(_1064_ | _0890_);
  assign _1067_ = _1066_ & ~(_0514_);
  assign _1068_ = _1067_ | _1062_;
  assign _1069_ = last_r[0] | ~(reqs_i[5]);
  assign _1070_ = _1069_ | _0273_;
  assign _1071_ = _1120_ & ~(_1070_);
  assign _1072_ = _0390_ & ~(_1036_);
  assign _1073_ = _1072_ | _1071_;
  assign _1074_ = _1073_ | _1068_;
  assign _1075_ = _1074_ | _1058_;
  assign _1077_ = ~(_1069_ | _0308_);
  assign _1078_ = _1077_ & ~(_0462_);
  assign _1079_ = _1035_ | _0758_;
  assign _1080_ = _0528_ & ~(_1079_);
  assign _1081_ = _1080_ | _1078_;
  assign _1082_ = _1069_ | _1131_;
  assign _1083_ = _1082_ | _0405_;
  assign _1084_ = _1120_ & ~(_1083_);
  assign _1085_ = _1035_ | _0491_;
  assign _1086_ = _1085_ | _0769_;
  assign _1088_ = _0490_ & ~(_1086_);
  assign _1089_ = _1088_ | _1084_;
  assign _1090_ = _1089_ | _1081_;
  assign _1091_ = ~_0538_;
  assign _1092_ = _1035_ | _0868_;
  assign _1093_ = _1092_ | _0769_;
  assign _1094_ = _1091_ & ~(_1093_);
  assign _1095_ = _1035_ | _1076_;
  assign _1096_ = _0427_ & ~(_1095_);
  assign _1097_ = _0787_ | _1120_;
  assign _1099_ = _1096_ & ~(_1097_);
  assign _1100_ = _1099_ | _1094_;
  assign _1101_ = _1035_ | _0857_;
  assign _1102_ = _0427_ & ~(_1101_);
  assign _1103_ = _0794_ | _1010_;
  assign _1104_ = _1102_ & ~(_1103_);
  assign _1105_ = _1035_ | _1054_;
  assign _1106_ = _0427_ & ~(_1105_);
  assign _1107_ = _0659_ | _0478_;
  assign _1108_ = _1106_ & ~(_1107_);
  assign _1110_ = _1108_ | _1104_;
  assign _1111_ = _1110_ | _1100_;
  assign _1112_ = _1111_ | _1090_;
  assign _1113_ = _1112_ | _1075_;
  assign _1114_ = ~(reqs_i[4] & last_r[0]);
  assign _1115_ = _1114_ | _0922_;
  assign _1116_ = _1115_ | _0769_;
  assign _1117_ = last_r[3] & ~(_1116_);
  assign _1118_ = reqs_i[10] | ~(reqs_i[4]);
  assign _1119_ = _1118_ | _1054_;
  assign _1121_ = _0427_ & ~(_1119_);
  assign _1122_ = _1142_ | _1098_;
  assign _1123_ = _1121_ & ~(_1122_);
  assign _1124_ = _1123_ | _1117_;
  assign _1125_ = reqs_i[9] | ~(reqs_i[4]);
  assign _1126_ = _1125_ | _0835_;
  assign _1127_ = _0427_ & ~(_1126_);
  assign _1128_ = _0021_ | _0879_;
  assign _1129_ = _1127_ & ~(_1128_);
  assign _1130_ = reqs_i[8] | ~(reqs_i[4]);
  assign _1132_ = _1130_ | _0076_;
  assign _1133_ = _1132_ | _0769_;
  assign _1134_ = _0120_ | _0098_;
  assign _1135_ = _1134_ | _1133_;
  assign _1136_ = _1120_ & ~(_1135_);
  assign _1137_ = _1136_ | _1129_;
  assign _1138_ = _1137_ | _1124_;
  assign _1139_ = reqs_i[7] | ~(reqs_i[4]);
  assign _1140_ = _1139_ | _0824_;
  assign _1141_ = _1140_ | _0769_;
  assign _1143_ = _1141_ | _0302_;
  assign _1144_ = _0369_ & ~(_1143_);
  assign _1145_ = reqs_i[6] | ~(reqs_i[4]);
  assign _1146_ = _1145_ | _0252_;
  assign _1147_ = _1146_ | _0769_;
  assign _1148_ = _1147_ | _0312_;
  assign _1149_ = _0566_ & ~(_1148_);
  assign _1150_ = _1149_ | _1144_;
  assign _1151_ = reqs_i[5] | ~(reqs_i[4]);
  assign _1152_ = _1151_ | _0791_;
  assign _1154_ = _1152_ | _0769_;
  assign _1155_ = _1154_ | _0890_;
  assign _1156_ = _0282_ & ~(_1155_);
  assign _1157_ = _1114_ | _0293_;
  assign _1158_ = _1120_ & ~(_1157_);
  assign _1159_ = _1158_ | _1156_;
  assign _1160_ = _1159_ | _1150_;
  assign _1161_ = _1160_ | _1138_;
  assign _1162_ = reqs_i[3] | ~(reqs_i[4]);
  assign _1163_ = _1162_ | _0977_;
  assign _1165_ = _0390_ & ~(_1163_);
  assign _1166_ = ~(_1114_ | _0758_);
  assign _1167_ = _1166_ & ~(_0314_);
  assign _1168_ = _1167_ | _1165_;
  assign _1169_ = ~(_1162_ | _0404_);
  assign _1170_ = _1169_ & ~(_0320_);
  assign _1171_ = reqs_i[15] | ~(reqs_i[4]);
  assign _1172_ = _1171_ | _0977_;
  assign _1173_ = _1172_ | _0769_;
  assign _1174_ = _0587_ & ~(_1173_);
  assign _1176_ = _1174_ | _1170_;
  assign _1177_ = _1176_ | _1168_;
  assign _1178_ = reqs_i[14] | ~(reqs_i[4]);
  assign _1179_ = _1178_ | _1087_;
  assign _1180_ = _1179_ | _0769_;
  assign _1181_ = _0593_ & ~(_1180_);
  assign _1182_ = reqs_i[13] | ~(reqs_i[4]);
  assign _1183_ = _1182_ | _0868_;
  assign _1184_ = _1183_ | _0769_;
  assign _1185_ = _0600_ & ~(_1184_);
  assign _0000_ = _1185_ | _1181_;
  assign _0001_ = reqs_i[12] | ~(reqs_i[4]);
  assign _0002_ = _0001_ | _1076_;
  assign _0003_ = _0427_ & ~(_0002_);
  assign _0004_ = _0294_ | _1120_;
  assign _0005_ = _0003_ & ~(_0004_);
  assign _0006_ = reqs_i[11] | ~(reqs_i[4]);
  assign _0007_ = _0006_ | _0857_;
  assign _0008_ = _0427_ & ~(_0007_);
  assign _0009_ = _1010_ | _0988_;
  assign _0011_ = _0008_ & ~(_0009_);
  assign _0012_ = _0011_ | _0005_;
  assign _0013_ = _0012_ | _0000_;
  assign _0014_ = _0013_ | _1177_;
  assign _0015_ = _0014_ | _1161_;
  assign _0016_ = _0015_ | _1113_;
  assign _0017_ = _0016_ | _1034_;
  assign _0018_ = reqs_i[2] | ~(reqs_i[3]);
  assign _0019_ = _0018_ | _0747_;
  assign _0020_ = ~(_0019_ | _0351_);
  assign _0022_ = _0378_ & ~(_0019_);
  assign _0023_ = _0654_ | _1010_;
  assign _0024_ = _0022_ & ~(_0023_);
  assign _0025_ = _0024_ | _0020_;
  assign _0026_ = _0382_ & ~(_0019_);
  assign _0027_ = _0659_ | _1142_;
  assign _0028_ = _0026_ & ~(_0027_);
  assign _0029_ = _0277_ & ~(_0019_);
  assign _0030_ = _0370_ | _0879_;
  assign _0031_ = _0029_ & ~(_0030_);
  assign _0033_ = _0031_ | _0028_;
  assign _0034_ = _0033_ | _0025_;
  assign _0035_ = _0019_ | _0291_;
  assign _0036_ = _0650_ | _0098_;
  assign _0037_ = _0036_ | _0035_;
  assign _0038_ = _1120_ & ~(_0037_);
  assign _0039_ = _0019_ | _0300_;
  assign _0040_ = _0039_ | _0891_;
  assign _0041_ = _0369_ & ~(_0040_);
  assign _0042_ = _0041_ | _0038_;
  assign _0044_ = _0019_ | _0310_;
  assign _0045_ = _0044_ | _0895_;
  assign _0046_ = _0566_ & ~(_0045_);
  assign _0047_ = _0019_ | _0802_;
  assign _0048_ = _0047_ | _0890_;
  assign _0049_ = _0391_ & ~(_0048_);
  assign _0050_ = _0049_ | _0046_;
  assign _0051_ = _0050_ | _0042_;
  assign _0052_ = _0051_ | _0034_;
  assign _0053_ = last_r[0] | ~(reqs_i[3]);
  assign _0055_ = _0053_ | _0293_;
  assign _0056_ = _1120_ & ~(_0055_);
  assign _0057_ = _0018_ | _0359_;
  assign _0058_ = _0390_ & ~(_0057_);
  assign _0059_ = _0058_ | _0056_;
  assign _0060_ = ~(_0053_ | _0404_);
  assign _0061_ = _0060_ & ~(_0314_);
  assign _0062_ = _0019_ | _0650_;
  assign _0063_ = last_r[3] & ~(_0062_);
  assign _0064_ = _0063_ | _0061_;
  assign _0066_ = _0064_ | _0059_;
  assign _0067_ = _0019_ | _0654_;
  assign _0068_ = ~(_0067_ | _0327_);
  assign _0069_ = _0019_ | _0659_;
  assign _0070_ = _0593_ & ~(_0069_);
  assign _0071_ = _0070_ | _0068_;
  assign _0072_ = _0019_ | _0879_;
  assign _0073_ = _0415_ & ~(_0072_);
  assign _0074_ = _0372_ & ~(_0019_);
  assign _0075_ = _0937_ | _1120_;
  assign _0077_ = _0074_ & ~(_0075_);
  assign _0078_ = _0077_ | _0073_;
  assign _0079_ = _0078_ | _0071_;
  assign _0080_ = _0079_ | _0066_;
  assign _0081_ = _0080_ | _0052_;
  assign _0082_ = ~(reqs_i[2] & last_r[0]);
  assign _0083_ = _0082_ | _0747_;
  assign _0084_ = ~(_0083_ | _0425_);
  assign _0085_ = reqs_i[10] | ~(reqs_i[2]);
  assign _0086_ = _0085_ | _0747_;
  assign _0088_ = _0372_ & ~(_0086_);
  assign _0089_ = _0953_ | _1120_;
  assign _0090_ = _0088_ & ~(_0089_);
  assign _0091_ = _0090_ | _0084_;
  assign _0092_ = reqs_i[9] | ~(reqs_i[2]);
  assign _0093_ = _0092_ | _0747_;
  assign _0094_ = _0378_ & ~(_0093_);
  assign _0095_ = _0718_ | _1010_;
  assign _0096_ = _0094_ & ~(_0095_);
  assign _0097_ = reqs_i[8] | ~(reqs_i[2]);
  assign _0099_ = _0097_ | _0747_;
  assign _0100_ = _0382_ & ~(_0099_);
  assign _0101_ = _0448_ | _1098_;
  assign _0102_ = _0100_ & ~(_0101_);
  assign _0103_ = _0102_ | _0096_;
  assign _0104_ = _0103_ | _0091_;
  assign _0105_ = reqs_i[7] | ~(reqs_i[2]);
  assign _0106_ = _0105_ | _0747_;
  assign _0107_ = _0277_ & ~(_0106_);
  assign _0108_ = _0452_ | _0879_;
  assign _0110_ = _0107_ & ~(_0108_);
  assign _0111_ = reqs_i[6] | ~(reqs_i[2]);
  assign _0112_ = _0111_ | _0747_;
  assign _0113_ = _0112_ | _0291_;
  assign _0114_ = _0712_ | _0098_;
  assign _0115_ = _0114_ | _0113_;
  assign _0116_ = _1120_ & ~(_0115_);
  assign _0117_ = _0116_ | _0110_;
  assign _0118_ = reqs_i[5] | ~(reqs_i[2]);
  assign _0119_ = _0118_ | _0747_;
  assign _0121_ = _0119_ | _0300_;
  assign _0122_ = _0121_ | _0962_;
  assign _0123_ = _0369_ & ~(_0122_);
  assign _0124_ = reqs_i[4] | ~(reqs_i[2]);
  assign _0125_ = _0124_ | _0747_;
  assign _0126_ = _0125_ | _0310_;
  assign _0127_ = _0126_ | _0312_;
  assign _0128_ = _0691_ & ~(_0127_);
  assign _0129_ = _0128_ | _0123_;
  assign _0130_ = _0129_ | _0117_;
  assign _0132_ = _0130_ | _0104_;
  assign _0133_ = reqs_i[3] | ~(reqs_i[2]);
  assign _0134_ = _0133_ | _0747_;
  assign _0135_ = _0134_ | _0802_;
  assign _0136_ = _0135_ | _0890_;
  assign _0137_ = _0466_ & ~(_0136_);
  assign _0138_ = _0082_ | _1131_;
  assign _0139_ = _1120_ & ~(_0138_);
  assign _0140_ = _0139_ | _0137_;
  assign _0141_ = reqs_i[1] | ~(reqs_i[2]);
  assign _0143_ = _0141_ | _0010_;
  assign _0144_ = _0390_ & ~(_0143_);
  assign _0145_ = reqs_i[15] | ~(reqs_i[2]);
  assign _0146_ = ~(_0145_ | _0747_);
  assign _0147_ = _0146_ & ~(_0433_);
  assign _0148_ = _0147_ | _0144_;
  assign _0149_ = _0148_ | _0140_;
  assign _0150_ = reqs_i[14] | ~(reqs_i[2]);
  assign _0151_ = _0150_ | _0747_;
  assign _0152_ = _0151_ | _0712_;
  assign _0154_ = last_r[3] & ~(_0152_);
  assign _0155_ = reqs_i[13] | ~(reqs_i[2]);
  assign _0156_ = _0155_ | _0747_;
  assign _0157_ = _0156_ | _0718_;
  assign _0158_ = _0587_ & ~(_0157_);
  assign _0159_ = _0158_ | _0154_;
  assign _0160_ = reqs_i[12] | ~(reqs_i[2]);
  assign _0161_ = _0160_ | _0747_;
  assign _0162_ = _0161_ | _1098_;
  assign _0163_ = _0723_ & ~(_0162_);
  assign _0165_ = reqs_i[11] | ~(reqs_i[2]);
  assign _0166_ = _0165_ | _0747_;
  assign _0167_ = _0166_ | _0879_;
  assign _0168_ = _0438_ & ~(_0167_);
  assign _0169_ = _0168_ | _0163_;
  assign _0170_ = _0169_ | _0159_;
  assign _0171_ = _0170_ | _0149_;
  assign _0172_ = _0171_ | _0132_;
  assign _0173_ = _0172_ | _0081_;
  assign _0174_ = reqs_i[0] | ~(reqs_i[1]);
  assign _0176_ = _0174_ | _0350_;
  assign _0177_ = ~(_0176_ | _0327_);
  assign _0178_ = _0174_ | _0835_;
  assign _0179_ = _0178_ | _0879_;
  assign _0180_ = _0501_ & ~(_0179_);
  assign _0181_ = _0180_ | _0177_;
  assign _0182_ = _0174_ | _0076_;
  assign _0183_ = _0372_ & ~(_0182_);
  assign _0184_ = _1047_ | _1120_;
  assign _0185_ = _0183_ & ~(_0184_);
  assign _0187_ = _0174_ | _0824_;
  assign _0188_ = _0378_ & ~(_0187_);
  assign _0189_ = _0794_ | _0197_;
  assign _0190_ = _0188_ & ~(_0189_);
  assign _0191_ = _0190_ | _0185_;
  assign _0192_ = _0191_ | _0181_;
  assign _0193_ = _0174_ | _0252_;
  assign _0194_ = _0382_ & ~(_0193_);
  assign _0195_ = _0659_ | _0448_;
  assign _0196_ = _0194_ & ~(_0195_);
  assign _0198_ = _0174_ | _0791_;
  assign _0199_ = _0277_ & ~(_0198_);
  assign _0200_ = _0514_ | _0879_;
  assign _0201_ = _0199_ & ~(_0200_);
  assign _0202_ = _0201_ | _0196_;
  assign _0203_ = _0174_ | _0289_;
  assign _0204_ = _0203_ | _0291_;
  assign _0205_ = _0787_ | _0098_;
  assign _0206_ = _0205_ | _0204_;
  assign _0207_ = _1120_ & ~(_0206_);
  assign _0209_ = _0174_ | _0780_;
  assign _0210_ = _0209_ | _0300_;
  assign _0211_ = _0210_ | _1053_;
  assign _0212_ = _0390_ & ~(_0211_);
  assign _0213_ = _0212_ | _0207_;
  assign _0214_ = _0213_ | _0202_;
  assign _0215_ = _0214_ | _0192_;
  assign _0216_ = _0174_ | _0308_;
  assign _0217_ = _0216_ | _0310_;
  assign _0218_ = _0217_ | _0895_;
  assign _0220_ = _0691_ & ~(_0218_);
  assign _0221_ = _0174_ | _0758_;
  assign _0222_ = _0221_ | _0802_;
  assign _0223_ = _0222_ | _0890_;
  assign _0224_ = _0528_ & ~(_0223_);
  assign _0225_ = _0224_ | _0220_;
  assign _0226_ = last_r[0] | ~(reqs_i[1]);
  assign _0227_ = _0226_ | _1131_;
  assign _0228_ = _1120_ & ~(_0227_);
  assign _0229_ = ~(_0174_ | _0491_);
  assign _0231_ = _0229_ & ~(_0425_);
  assign _0232_ = _0231_ | _0228_;
  assign _0233_ = _0232_ | _0225_;
  assign _0234_ = ~(_0174_ | _0868_);
  assign _0235_ = _0234_ & ~(_0538_);
  assign _0236_ = _0174_ | _1076_;
  assign _0237_ = _0236_ | _0787_;
  assign _0238_ = last_r[3] & ~(_0237_);
  assign _0239_ = _0238_ | _0235_;
  assign _0240_ = _0174_ | _0857_;
  assign _0242_ = _0240_ | _0794_;
  assign _0243_ = _0358_ & ~(_0242_);
  assign _0244_ = _0174_ | _1054_;
  assign _0245_ = _0244_ | _0659_;
  assign _0246_ = _0723_ & ~(_0245_);
  assign _0247_ = _0246_ | _0243_;
  assign _0248_ = _0247_ | _0239_;
  assign _0249_ = _0248_ | _0233_;
  assign _0250_ = _0249_ | _0215_;
  assign _0251_ = _0250_ | _0345_;
  assign _0253_ = _0251_ | _0173_;
  assign _0254_ = _0253_ | _0017_;
  assign _0255_ = _0885_ & ~(_0254_);
  assign sel_one_hot_o[0] = _0345_ & ~(_0255_);
  assign sel_one_hot_o[1] = _0250_ & ~(_0255_);
  assign sel_one_hot_o[2] = _0172_ & ~(_0255_);
  assign sel_one_hot_o[3] = _0081_ & ~(_0255_);
  assign sel_one_hot_o[4] = _0015_ & ~(_0255_);
  assign sel_one_hot_o[5] = _1113_ & ~(_0255_);
  assign sel_one_hot_o[6] = _1033_ & ~(_0255_);
  assign sel_one_hot_o[7] = _0945_ & ~(_0255_);
  assign sel_one_hot_o[8] = _0882_ & ~(_0255_);
  assign sel_one_hot_o[9] = _0806_ & ~(_0255_);
  assign sel_one_hot_o[10] = _0737_ & ~(_0255_);
  assign sel_one_hot_o[11] = _0669_ & ~(_0255_);
  assign sel_one_hot_o[12] = _0610_ & ~(_0255_);
  assign sel_one_hot_o[13] = _0546_ & ~(_0255_);
  assign sel_one_hot_o[14] = _0483_ & ~(_0255_);
  assign sel_one_hot_o[15] = _0420_ & ~(_0255_);
  assign _0257_ = _0546_ | _0420_;
  assign _0259_ = _0806_ | _0669_;
  assign _0260_ = _0259_ | _0257_;
  assign _0261_ = _1113_ | _0945_;
  assign _0262_ = _0250_ | _0081_;
  assign _0263_ = _0262_ | _0261_;
  assign _0264_ = _0263_ | _0260_;
  assign _0265_ = _0250_ | _0173_;
  assign _0266_ = _0265_ | _0017_;
  assign _0267_ = _0266_ | ~(_0885_);
  assign tag_o[0] = _0267_ & _0264_;
  assign _0269_ = _0484_ & ~(_0738_);
  assign _0270_ = _0173_ | _1034_;
  assign _0271_ = _0269_ & ~(_0270_);
  assign tag_o[1] = _0267_ & ~(_0271_);
  assign _0272_ = _0612_ & ~(_0017_);
  assign tag_o[2] = _0267_ & ~(_0272_);
  assign tag_o[3] = _0267_ & ~(_0885_);
  assign grants_o[0] = sel_one_hot_o[0] & grants_en_i;
  assign grants_o[1] = sel_one_hot_o[1] & grants_en_i;
  assign grants_o[2] = sel_one_hot_o[2] & grants_en_i;
  assign grants_o[3] = sel_one_hot_o[3] & grants_en_i;
  assign grants_o[4] = sel_one_hot_o[4] & grants_en_i;
  assign grants_o[5] = sel_one_hot_o[5] & grants_en_i;
  assign grants_o[6] = sel_one_hot_o[6] & grants_en_i;
  assign grants_o[7] = sel_one_hot_o[7] & grants_en_i;
  assign grants_o[8] = sel_one_hot_o[8] & grants_en_i;
  assign grants_o[9] = sel_one_hot_o[9] & grants_en_i;
  assign grants_o[10] = sel_one_hot_o[10] & grants_en_i;
  assign grants_o[11] = sel_one_hot_o[11] & grants_en_i;
  assign grants_o[12] = sel_one_hot_o[12] & grants_en_i;
  assign grants_o[13] = sel_one_hot_o[13] & grants_en_i;
  assign grants_o[14] = sel_one_hot_o[14] & grants_en_i;
  assign grants_o[15] = sel_one_hot_o[15] & grants_en_i;
  always @(posedge clk_i)
    if (reset_i) last_r[0] <= 1'h0;
    else if (yumi_i) last_r[0] <= tag_o[0];
  always @(posedge clk_i)
    if (reset_i) last_r[1] <= 1'h0;
    else if (yumi_i) last_r[1] <= tag_o[1];
  always @(posedge clk_i)
    if (reset_i) last_r[2] <= 1'h0;
    else if (yumi_i) last_r[2] <= tag_o[2];
  always @(posedge clk_i)
    if (reset_i) last_r[3] <= 1'h0;
    else if (yumi_i) last_r[3] <= tag_o[3];
  assign hold_on_sr = 1'h0;
  assign \inputs_16.sel_one_hot_n  = sel_one_hot_o;
  assign reset_on_sr = 1'h0;
endmodule
