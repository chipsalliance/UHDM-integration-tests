module bsg_tiehi(o);
  output [15:0] o;
  wire [15:0] o;
  assign o = 16'hffff;
endmodule
