module bsg_abs(a_i, o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  input [15:0] a_i;
  wire [15:0] a_i;
  output [15:0] o;
  wire [15:0] o;
  assign _00_ = a_i[0] ^ a_i[1];
  assign o[1] = a_i[15] ? _00_ : a_i[1];
  assign _01_ = a_i[0] | a_i[1];
  assign _02_ = _01_ ^ a_i[2];
  assign o[2] = a_i[15] ? _02_ : a_i[2];
  assign _03_ = _01_ | a_i[2];
  assign _04_ = _03_ ^ a_i[3];
  assign o[3] = a_i[15] ? _04_ : a_i[3];
  assign _05_ = a_i[3] | a_i[2];
  assign _06_ = _05_ | _01_;
  assign _07_ = _06_ ^ a_i[4];
  assign o[4] = a_i[15] ? _07_ : a_i[4];
  assign _08_ = _06_ | a_i[4];
  assign _09_ = _08_ ^ a_i[5];
  assign o[5] = a_i[15] ? _09_ : a_i[5];
  assign _10_ = a_i[5] | a_i[4];
  assign _11_ = _10_ | _06_;
  assign _12_ = _11_ ^ a_i[6];
  assign o[6] = a_i[15] ? _12_ : a_i[6];
  assign _13_ = _11_ | a_i[6];
  assign _14_ = _13_ ^ a_i[7];
  assign o[7] = a_i[15] ? _14_ : a_i[7];
  assign _15_ = a_i[7] | a_i[6];
  assign _16_ = _15_ | _10_;
  assign _17_ = _16_ | _06_;
  assign _18_ = _17_ ^ a_i[8];
  assign o[8] = a_i[15] ? _18_ : a_i[8];
  assign _19_ = _17_ | a_i[8];
  assign _20_ = _19_ ^ a_i[9];
  assign o[9] = a_i[15] ? _20_ : a_i[9];
  assign _21_ = a_i[9] | a_i[8];
  assign _22_ = _21_ | _17_;
  assign _23_ = _22_ ^ a_i[10];
  assign o[10] = a_i[15] ? _23_ : a_i[10];
  assign _24_ = _22_ | a_i[10];
  assign _25_ = _24_ ^ a_i[11];
  assign o[11] = a_i[15] ? _25_ : a_i[11];
  assign _26_ = a_i[11] | a_i[10];
  assign _27_ = _26_ | _21_;
  assign _28_ = _27_ | _17_;
  assign _29_ = _28_ ^ a_i[12];
  assign o[12] = a_i[15] ? _29_ : a_i[12];
  assign _30_ = _28_ | a_i[12];
  assign _31_ = _30_ ^ a_i[13];
  assign o[13] = a_i[15] ? _31_ : a_i[13];
  assign _32_ = a_i[13] | a_i[12];
  assign _33_ = _32_ | _28_;
  assign _34_ = _33_ ^ a_i[14];
  assign o[14] = a_i[15] ? _34_ : a_i[14];
  assign _35_ = _33_ | a_i[14];
  assign o[15] = a_i[15] & ~(_35_);
  assign o[0] = a_i[0];
endmodule
