module bsg_counter_up_down_variable(clk_i, reset_i, up_i, down_i, count_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire [9:0] _050_;
  wire [9:0] _051_;
  input clk_i;
  wire clk_i;
  output [9:0] count_o;
  reg [9:0] count_o;
  input down_i;
  wire down_i;
  input reset_i;
  wire reset_i;
  input up_i;
  wire up_i;
  assign _000_ = down_i & ~(up_i);
  assign _001_ = _000_ ^ count_o[1];
  assign _002_ = ~count_o[0];
  assign _003_ = ~(down_i ^ up_i);
  assign _004_ = _003_ | _002_;
  assign _051_[1] = ~(_004_ ^ _001_);
  assign _005_ = count_o[1] ^ count_o[2];
  assign _006_ = ~(_000_ | count_o[1]);
  assign _007_ = _001_ & ~(_004_);
  assign _008_ = _007_ | _006_;
  assign _051_[2] = ~(_008_ ^ _005_);
  assign _009_ = count_o[2] ^ count_o[3];
  assign _010_ = count_o[2] | ~(count_o[1]);
  assign _011_ = _008_ & ~(_005_);
  assign _012_ = _010_ & ~(_011_);
  assign _051_[3] = _012_ ^ _009_;
  assign _013_ = count_o[3] ^ count_o[4];
  assign _014_ = count_o[2] & ~(count_o[3]);
  assign _015_ = ~(_010_ | _009_);
  assign _016_ = ~(_015_ | _014_);
  assign _017_ = _009_ | _005_;
  assign _018_ = _008_ & ~(_017_);
  assign _019_ = _016_ & ~(_018_);
  assign _051_[4] = _019_ ^ _013_;
  assign _020_ = count_o[4] ^ count_o[5];
  assign _021_ = count_o[4] | ~(count_o[3]);
  assign _022_ = _018_ | ~(_016_);
  assign _023_ = _022_ & ~(_013_);
  assign _024_ = _021_ & ~(_023_);
  assign _051_[5] = _024_ ^ _020_;
  assign _025_ = count_o[5] ^ count_o[6];
  assign _026_ = count_o[4] & ~(count_o[5]);
  assign _027_ = ~(_021_ | _020_);
  assign _028_ = _027_ | _026_;
  assign _029_ = _020_ | _013_;
  assign _030_ = _029_ | _019_;
  assign _031_ = _030_ & ~(_028_);
  assign _051_[6] = _031_ ^ _025_;
  assign _032_ = count_o[6] ^ count_o[7];
  assign _033_ = count_o[6] | ~(count_o[5]);
  assign _034_ = ~(_031_ | _025_);
  assign _035_ = _033_ & ~(_034_);
  assign _051_[7] = _035_ ^ _032_;
  assign _036_ = count_o[8] ^ count_o[7];
  assign _037_ = count_o[7] | ~(count_o[6]);
  assign _038_ = ~(_033_ | _032_);
  assign _039_ = _037_ & ~(_038_);
  assign _040_ = _032_ | _025_;
  assign _041_ = _028_ & ~(_040_);
  assign _042_ = _039_ & ~(_041_);
  assign _043_ = _040_ | _029_;
  assign _044_ = _022_ & ~(_043_);
  assign _045_ = _042_ & ~(_044_);
  assign _051_[8] = _045_ ^ _036_;
  assign _046_ = count_o[9] ^ count_o[8];
  assign _047_ = count_o[8] | ~(count_o[7]);
  assign _048_ = ~(_045_ | _036_);
  assign _049_ = _047_ & ~(_048_);
  assign _051_[9] = _049_ ^ _046_;
  assign _050_[0] = _003_ ^ _002_;
  always @(posedge clk_i)
    if (reset_i) count_o[4] <= 1'h0;
    else count_o[4] <= _051_[4];
  always @(posedge clk_i)
    if (reset_i) count_o[5] <= 1'h0;
    else count_o[5] <= _051_[5];
  always @(posedge clk_i)
    if (reset_i) count_o[6] <= 1'h0;
    else count_o[6] <= _051_[6];
  always @(posedge clk_i)
    if (reset_i) count_o[7] <= 1'h0;
    else count_o[7] <= _051_[7];
  always @(posedge clk_i)
    if (reset_i) count_o[8] <= 1'h0;
    else count_o[8] <= _051_[8];
  always @(posedge clk_i)
    if (reset_i) count_o[9] <= 1'h0;
    else count_o[9] <= _051_[9];
  always @(posedge clk_i)
    if (reset_i) count_o[0] <= 1'h0;
    else count_o[0] <= _050_[0];
  always @(posedge clk_i)
    if (reset_i) count_o[1] <= 1'h0;
    else count_o[1] <= _051_[1];
  always @(posedge clk_i)
    if (reset_i) count_o[2] <= 1'h0;
    else count_o[2] <= _051_[2];
  always @(posedge clk_i)
    if (reset_i) count_o[3] <= 1'h0;
    else count_o[3] <= _051_[3];
  assign _051_[0] = _050_[0];
endmodule
