module bsg_make_2D_array(i, o);
  input [159:0] i;
  wire [159:0] i;
  output [159:0] o;
  wire [159:0] o;
  assign o = i;
endmodule
