module bsg_counter_overflow_set_en(clk_i, en_i, set_i, val_i, count_o, overflow_o);
  wire [23:0] _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  input clk_i;
  wire clk_i;
  output [23:0] count_o;
  reg [23:0] count_o;
  input en_i;
  wire en_i;
  output overflow_o;
  wire overflow_o;
  input set_i;
  wire set_i;
  input [23:0] val_i;
  wire [23:0] val_i;
  assign _091_ = count_o[1] | count_o[0];
  assign _092_ = count_o[3] | count_o[2];
  assign _093_ = _092_ | _091_;
  assign _094_ = count_o[5] | count_o[4];
  assign _095_ = count_o[6] | ~(count_o[7]);
  assign _096_ = _095_ | _094_;
  assign _097_ = _096_ | _093_;
  assign _098_ = count_o[8] | ~(count_o[9]);
  assign _099_ = count_o[11] | ~(count_o[10]);
  assign _100_ = _099_ | _098_;
  assign _101_ = count_o[13] | ~(count_o[12]);
  assign _102_ = count_o[14] | ~(count_o[15]);
  assign _103_ = _102_ | _101_;
  assign _104_ = _103_ | _100_;
  assign _105_ = _104_ | _097_;
  assign _106_ = count_o[17] | count_o[16];
  assign _107_ = count_o[18] | ~(count_o[19]);
  assign _108_ = _107_ | _106_;
  assign _109_ = count_o[21] | ~(count_o[20]);
  assign _110_ = count_o[22] | ~(count_o[23]);
  assign _111_ = _110_ | _109_;
  assign _112_ = _111_ | _108_;
  assign _113_ = _112_ | _105_;
  assign overflow_o = ~_113_;
  assign _002_ = set_i | en_i;
  assign _001_ = _002_ | ~(_113_);
  assign _003_ = _113_ & ~(count_o[0]);
  assign _000_[0] = set_i ? val_i[0] : _003_;
  assign _004_ = ~(count_o[1] ^ count_o[0]);
  assign _005_ = _113_ & ~(_004_);
  assign _000_[1] = set_i ? val_i[1] : _005_;
  assign _006_ = ~(count_o[1] & count_o[0]);
  assign _007_ = _006_ ^ count_o[2];
  assign _008_ = _113_ & ~(_007_);
  assign _000_[2] = set_i ? val_i[2] : _008_;
  assign _009_ = count_o[1] & count_o[0];
  assign _010_ = ~(_009_ & count_o[2]);
  assign _011_ = _010_ ^ count_o[3];
  assign _012_ = _113_ & ~(_011_);
  assign _000_[3] = set_i ? val_i[3] : _012_;
  assign _013_ = ~(count_o[3] & count_o[2]);
  assign _014_ = _013_ | _006_;
  assign _015_ = _014_ ^ count_o[4];
  assign _016_ = _113_ & ~(_015_);
  assign _000_[4] = set_i ? val_i[4] : _016_;
  assign _017_ = _009_ & ~(_013_);
  assign _018_ = ~(_017_ & count_o[4]);
  assign _019_ = _018_ ^ count_o[5];
  assign _020_ = _113_ & ~(_019_);
  assign _000_[5] = set_i ? val_i[5] : _020_;
  assign _021_ = ~(count_o[5] & count_o[4]);
  assign _022_ = _021_ | _014_;
  assign _023_ = _022_ ^ count_o[6];
  assign _024_ = _113_ & ~(_023_);
  assign _000_[6] = set_i ? val_i[6] : _024_;
  assign _025_ = _022_ | ~(count_o[6]);
  assign _026_ = _025_ ^ count_o[7];
  assign _027_ = _113_ & ~(_026_);
  assign _000_[7] = set_i ? val_i[7] : _027_;
  assign _028_ = ~(count_o[7] & count_o[6]);
  assign _029_ = _028_ | _021_;
  assign _030_ = _029_ | _014_;
  assign _031_ = _030_ ^ count_o[8];
  assign _032_ = _113_ & ~(_031_);
  assign _000_[8] = set_i ? val_i[8] : _032_;
  assign _033_ = _017_ & ~(_029_);
  assign _034_ = ~(_033_ & count_o[8]);
  assign _035_ = _034_ ^ count_o[9];
  assign _036_ = _113_ & ~(_035_);
  assign _000_[9] = set_i ? val_i[9] : _036_;
  assign _037_ = ~(count_o[9] & count_o[8]);
  assign _038_ = _037_ | _030_;
  assign _039_ = _038_ ^ count_o[10];
  assign _040_ = _113_ & ~(_039_);
  assign _000_[10] = set_i ? val_i[10] : _040_;
  assign _041_ = _038_ | ~(count_o[10]);
  assign _042_ = _041_ ^ count_o[11];
  assign _043_ = _113_ & ~(_042_);
  assign _000_[11] = set_i ? val_i[11] : _043_;
  assign _044_ = ~(count_o[11] & count_o[10]);
  assign _045_ = _044_ | _037_;
  assign _046_ = _045_ | _030_;
  assign _047_ = _046_ ^ count_o[12];
  assign _048_ = _113_ & ~(_047_);
  assign _000_[12] = set_i ? val_i[12] : _048_;
  assign _049_ = _046_ | ~(count_o[12]);
  assign _050_ = _049_ ^ count_o[13];
  assign _051_ = _113_ & ~(_050_);
  assign _000_[13] = set_i ? val_i[13] : _051_;
  assign _052_ = ~(count_o[13] & count_o[12]);
  assign _053_ = _052_ | _046_;
  assign _054_ = _053_ ^ count_o[14];
  assign _055_ = _113_ & ~(_054_);
  assign _000_[14] = set_i ? val_i[14] : _055_;
  assign _056_ = _053_ | ~(count_o[14]);
  assign _057_ = _056_ ^ count_o[15];
  assign _058_ = _113_ & ~(_057_);
  assign _000_[15] = set_i ? val_i[15] : _058_;
  assign _059_ = ~(count_o[14] & count_o[15]);
  assign _060_ = _059_ | _052_;
  assign _061_ = _060_ | _045_;
  assign _062_ = _061_ | _030_;
  assign _063_ = _062_ ^ count_o[16];
  assign _064_ = _113_ & ~(_063_);
  assign _000_[16] = set_i ? val_i[16] : _064_;
  assign _065_ = _033_ & ~(_061_);
  assign _066_ = ~(_065_ & count_o[16]);
  assign _067_ = _066_ ^ count_o[17];
  assign _068_ = _113_ & ~(_067_);
  assign _000_[17] = set_i ? val_i[17] : _068_;
  assign _069_ = ~(count_o[17] & count_o[16]);
  assign _070_ = _069_ | _062_;
  assign _071_ = _070_ ^ count_o[18];
  assign _072_ = _113_ & ~(_071_);
  assign _000_[18] = set_i ? val_i[18] : _072_;
  assign _073_ = _070_ | ~(count_o[18]);
  assign _074_ = _073_ ^ count_o[19];
  assign _075_ = _113_ & ~(_074_);
  assign _000_[19] = set_i ? val_i[19] : _075_;
  assign _076_ = ~(count_o[19] & count_o[18]);
  assign _077_ = _076_ | _069_;
  assign _078_ = _077_ | _062_;
  assign _079_ = _078_ ^ count_o[20];
  assign _080_ = _113_ & ~(_079_);
  assign _000_[20] = set_i ? val_i[20] : _080_;
  assign _081_ = _078_ | ~(count_o[20]);
  assign _082_ = _081_ ^ count_o[21];
  assign _083_ = _113_ & ~(_082_);
  assign _000_[21] = set_i ? val_i[21] : _083_;
  assign _084_ = ~(count_o[21] & count_o[20]);
  assign _085_ = _084_ | _078_;
  assign _086_ = _085_ ^ count_o[22];
  assign _087_ = _113_ & ~(_086_);
  assign _000_[22] = set_i ? val_i[22] : _087_;
  assign _088_ = _085_ | ~(count_o[22]);
  assign _089_ = _088_ ^ count_o[23];
  assign _090_ = _113_ & ~(_089_);
  assign _000_[23] = set_i ? val_i[23] : _090_;
  always @(posedge clk_i)
    if (_001_) count_o[0] <= _000_[0];
  always @(posedge clk_i)
    if (_001_) count_o[1] <= _000_[1];
  always @(posedge clk_i)
    if (_001_) count_o[2] <= _000_[2];
  always @(posedge clk_i)
    if (_001_) count_o[3] <= _000_[3];
  always @(posedge clk_i)
    if (_001_) count_o[4] <= _000_[4];
  always @(posedge clk_i)
    if (_001_) count_o[5] <= _000_[5];
  always @(posedge clk_i)
    if (_001_) count_o[6] <= _000_[6];
  always @(posedge clk_i)
    if (_001_) count_o[7] <= _000_[7];
  always @(posedge clk_i)
    if (_001_) count_o[8] <= _000_[8];
  always @(posedge clk_i)
    if (_001_) count_o[9] <= _000_[9];
  always @(posedge clk_i)
    if (_001_) count_o[10] <= _000_[10];
  always @(posedge clk_i)
    if (_001_) count_o[11] <= _000_[11];
  always @(posedge clk_i)
    if (_001_) count_o[12] <= _000_[12];
  always @(posedge clk_i)
    if (_001_) count_o[13] <= _000_[13];
  always @(posedge clk_i)
    if (_001_) count_o[14] <= _000_[14];
  always @(posedge clk_i)
    if (_001_) count_o[15] <= _000_[15];
  always @(posedge clk_i)
    if (_001_) count_o[16] <= _000_[16];
  always @(posedge clk_i)
    if (_001_) count_o[17] <= _000_[17];
  always @(posedge clk_i)
    if (_001_) count_o[18] <= _000_[18];
  always @(posedge clk_i)
    if (_001_) count_o[19] <= _000_[19];
  always @(posedge clk_i)
    if (_001_) count_o[20] <= _000_[20];
  always @(posedge clk_i)
    if (_001_) count_o[21] <= _000_[21];
  always @(posedge clk_i)
    if (_001_) count_o[22] <= _000_[22];
  always @(posedge clk_i)
    if (_001_) count_o[23] <= _000_[23];
endmodule
