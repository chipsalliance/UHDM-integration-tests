// We are actually testing including duplicated packages in Makefile,
// not this module
module top;
endmodule
