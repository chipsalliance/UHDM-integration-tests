module bsg_counter_dynamic_limit_en(clk_i, reset_i, en_i, limit_i, counter_o, overflowed_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  input clk_i;
  wire clk_i;
  output [15:0] counter_o;
  reg [15:0] counter_o;
  input en_i;
  wire en_i;
  input [15:0] limit_i;
  wire [15:0] limit_i;
  output overflowed_o;
  wire overflowed_o;
  input reset_i;
  wire reset_i;
  assign _021_ = limit_i[0] ^ counter_o[0];
  assign _022_ = ~(counter_o[1] ^ counter_o[0]);
  assign _023_ = ~(_022_ ^ limit_i[1]);
  assign _024_ = _021_ & ~(_023_);
  assign _025_ = ~(counter_o[1] & counter_o[0]);
  assign _026_ = _025_ ^ counter_o[2];
  assign _027_ = ~(_026_ ^ limit_i[2]);
  assign _028_ = counter_o[2] & ~(_025_);
  assign _029_ = ~(_028_ ^ counter_o[3]);
  assign _030_ = ~(_029_ ^ limit_i[3]);
  assign _031_ = _030_ | _027_;
  assign _032_ = _024_ & ~(_031_);
  assign _033_ = ~counter_o[4];
  assign _034_ = counter_o[3] & counter_o[2];
  assign _035_ = _034_ & ~(_025_);
  assign _036_ = _035_ ^ _033_;
  assign _037_ = ~(_036_ ^ limit_i[4]);
  assign _038_ = _035_ & ~(_033_);
  assign _039_ = ~(_038_ ^ counter_o[5]);
  assign _040_ = ~(_039_ ^ limit_i[5]);
  assign _041_ = _040_ | _037_;
  assign _042_ = ~(counter_o[5] & counter_o[4]);
  assign _043_ = _042_ | ~(_035_);
  assign _044_ = _043_ ^ counter_o[6];
  assign _045_ = ~(_044_ ^ limit_i[6]);
  assign _046_ = counter_o[6] & ~(_043_);
  assign _047_ = ~(_046_ ^ counter_o[7]);
  assign _048_ = ~(_047_ ^ limit_i[7]);
  assign _049_ = _048_ | _045_;
  assign _050_ = _049_ | _041_;
  assign _051_ = _032_ & ~(_050_);
  assign _052_ = ~counter_o[8];
  assign _053_ = ~(counter_o[7] & counter_o[6]);
  assign _054_ = _053_ | _042_;
  assign _055_ = _035_ & ~(_054_);
  assign _056_ = _055_ ^ _052_;
  assign _057_ = ~(_056_ ^ limit_i[8]);
  assign _058_ = _055_ & ~(_052_);
  assign _059_ = ~(_058_ ^ counter_o[9]);
  assign _060_ = ~(_059_ ^ limit_i[9]);
  assign _061_ = _060_ | _057_;
  assign _062_ = ~(counter_o[9] & counter_o[8]);
  assign _063_ = _062_ | ~(_055_);
  assign _064_ = _063_ ^ counter_o[10];
  assign _065_ = ~(_064_ ^ limit_i[10]);
  assign _066_ = counter_o[10] & ~(_063_);
  assign _067_ = ~(_066_ ^ counter_o[11]);
  assign _068_ = ~(_067_ ^ limit_i[11]);
  assign _069_ = _068_ | _065_;
  assign _070_ = _069_ | _061_;
  assign _000_ = ~counter_o[12];
  assign _001_ = ~(counter_o[11] & counter_o[10]);
  assign _002_ = _001_ | _062_;
  assign _003_ = _055_ & ~(_002_);
  assign _004_ = _003_ ^ _000_;
  assign _005_ = ~(_004_ ^ limit_i[12]);
  assign _006_ = _003_ & ~(_000_);
  assign _007_ = ~(_006_ ^ counter_o[13]);
  assign _008_ = ~(_007_ ^ limit_i[13]);
  assign _009_ = _008_ | _005_;
  assign _010_ = ~counter_o[14];
  assign _011_ = ~(counter_o[13] & counter_o[12]);
  assign _012_ = _003_ & ~(_011_);
  assign _013_ = _012_ ^ _010_;
  assign _014_ = ~(_013_ ^ limit_i[14]);
  assign _015_ = _012_ & ~(_010_);
  assign _016_ = ~(_015_ ^ counter_o[15]);
  assign _017_ = ~(_016_ ^ limit_i[15]);
  assign _018_ = _017_ | _014_;
  assign _019_ = _018_ | _009_;
  assign _020_ = _019_ | _070_;
  assign overflowed_o = _051_ & ~(_020_);
  assign _071_ = ~(overflowed_o | counter_o[0]);
  assign _078_ = ~(overflowed_o | _022_);
  assign _079_ = ~(overflowed_o | _026_);
  assign _080_ = ~(overflowed_o | _029_);
  assign _081_ = ~(overflowed_o | _036_);
  assign _082_ = ~(overflowed_o | _039_);
  assign _083_ = ~(overflowed_o | _044_);
  assign _084_ = ~(overflowed_o | _047_);
  assign _085_ = ~(overflowed_o | _056_);
  assign _086_ = ~(overflowed_o | _059_);
  assign _072_ = ~(overflowed_o | _064_);
  assign _073_ = ~(overflowed_o | _067_);
  assign _074_ = ~(overflowed_o | _004_);
  assign _075_ = ~(overflowed_o | _007_);
  assign _076_ = ~(overflowed_o | _013_);
  assign _077_ = ~(overflowed_o | _016_);
  always @(posedge clk_i)
    if (reset_i) counter_o[0] <= 1'h0;
    else if (en_i) counter_o[0] <= _071_;
  always @(posedge clk_i)
    if (reset_i) counter_o[1] <= 1'h0;
    else if (en_i) counter_o[1] <= _078_;
  always @(posedge clk_i)
    if (reset_i) counter_o[2] <= 1'h0;
    else if (en_i) counter_o[2] <= _079_;
  always @(posedge clk_i)
    if (reset_i) counter_o[3] <= 1'h0;
    else if (en_i) counter_o[3] <= _080_;
  always @(posedge clk_i)
    if (reset_i) counter_o[4] <= 1'h0;
    else if (en_i) counter_o[4] <= _081_;
  always @(posedge clk_i)
    if (reset_i) counter_o[5] <= 1'h0;
    else if (en_i) counter_o[5] <= _082_;
  always @(posedge clk_i)
    if (reset_i) counter_o[6] <= 1'h0;
    else if (en_i) counter_o[6] <= _083_;
  always @(posedge clk_i)
    if (reset_i) counter_o[7] <= 1'h0;
    else if (en_i) counter_o[7] <= _084_;
  always @(posedge clk_i)
    if (reset_i) counter_o[8] <= 1'h0;
    else if (en_i) counter_o[8] <= _085_;
  always @(posedge clk_i)
    if (reset_i) counter_o[9] <= 1'h0;
    else if (en_i) counter_o[9] <= _086_;
  always @(posedge clk_i)
    if (reset_i) counter_o[10] <= 1'h0;
    else if (en_i) counter_o[10] <= _072_;
  always @(posedge clk_i)
    if (reset_i) counter_o[11] <= 1'h0;
    else if (en_i) counter_o[11] <= _073_;
  always @(posedge clk_i)
    if (reset_i) counter_o[12] <= 1'h0;
    else if (en_i) counter_o[12] <= _074_;
  always @(posedge clk_i)
    if (reset_i) counter_o[13] <= 1'h0;
    else if (en_i) counter_o[13] <= _075_;
  always @(posedge clk_i)
    if (reset_i) counter_o[14] <= 1'h0;
    else if (en_i) counter_o[14] <= _076_;
  always @(posedge clk_i)
    if (reset_i) counter_o[15] <= 1'h0;
    else if (en_i) counter_o[15] <= _077_;
endmodule
