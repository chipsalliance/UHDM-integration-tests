module bsg_gray_to_binary(gray_i, binary_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  output [15:0] binary_o;
  wire [15:0] binary_o;
  input [15:0] gray_i;
  wire [15:0] gray_i;
  wire [15:0] \scan_xor.i ;
  wire [15:0] \scan_xor.o ;
  wire [15:0] \scan_xor.scanN.row[0].fill ;
  wire [15:0] \scan_xor.scanN.row[0].shifted ;
  wire [15:0] \scan_xor.scanN.row[1].fill ;
  wire [15:0] \scan_xor.scanN.row[1].shifted ;
  wire [15:0] \scan_xor.scanN.row[2].fill ;
  wire [15:0] \scan_xor.scanN.row[2].shifted ;
  wire [15:0] \scan_xor.scanN.row[3].fill ;
  wire [15:0] \scan_xor.scanN.row[3].shifted ;
  wire [79:0] \scan_xor.t ;
  assign _00_ = gray_i[13] ^ gray_i[12];
  assign _01_ = ~(gray_i[14] ^ gray_i[15]);
  assign _02_ = _01_ ^ _00_;
  assign binary_o[12] = ~_02_;
  assign _03_ = gray_i[9] ^ gray_i[8];
  assign _04_ = ~(gray_i[11] ^ gray_i[10]);
  assign _05_ = _04_ ^ _03_;
  assign binary_o[8] = _05_ ^ _02_;
  assign _06_ = ~(gray_i[14] ^ gray_i[13]);
  assign _07_ = _06_ ^ gray_i[15];
  assign binary_o[13] = ~_07_;
  assign _08_ = gray_i[10] ^ gray_i[9];
  assign _09_ = ~(gray_i[12] ^ gray_i[11]);
  assign _10_ = _09_ ^ _08_;
  assign binary_o[9] = _10_ ^ _07_;
  assign binary_o[14] = ~_01_;
  assign _11_ = _04_ ^ _00_;
  assign binary_o[10] = _11_ ^ _01_;
  assign _12_ = ~gray_i[15];
  assign _13_ = ~(_09_ ^ _06_);
  assign binary_o[11] = _13_ ^ _12_;
  assign _14_ = ~(gray_i[1] ^ gray_i[0]);
  assign _15_ = ~(gray_i[3] ^ gray_i[2]);
  assign _16_ = _15_ ^ _14_;
  assign _17_ = ~(gray_i[5] ^ gray_i[4]);
  assign _18_ = ~(gray_i[7] ^ gray_i[6]);
  assign _19_ = ~(_18_ ^ _17_);
  assign _20_ = ~(_19_ ^ _16_);
  assign binary_o[0] = _20_ ^ binary_o[8];
  assign _21_ = ~(gray_i[2] ^ gray_i[1]);
  assign _22_ = ~(gray_i[4] ^ gray_i[3]);
  assign _23_ = _22_ ^ _21_;
  assign _24_ = ~(gray_i[6] ^ gray_i[5]);
  assign _25_ = ~(gray_i[8] ^ gray_i[7]);
  assign _26_ = ~(_25_ ^ _24_);
  assign _27_ = ~(_26_ ^ _23_);
  assign binary_o[1] = _27_ ^ binary_o[9];
  assign _28_ = _17_ ^ _15_;
  assign _29_ = _18_ ^ _03_;
  assign _30_ = ~(_29_ ^ _28_);
  assign binary_o[2] = _30_ ^ binary_o[10];
  assign _31_ = _24_ ^ _22_;
  assign _32_ = _25_ ^ _08_;
  assign _33_ = ~(_32_ ^ _31_);
  assign binary_o[3] = _33_ ^ binary_o[11];
  assign _34_ = ~(_19_ ^ _05_);
  assign binary_o[4] = _34_ ^ _02_;
  assign _35_ = ~(_26_ ^ _10_);
  assign binary_o[5] = _35_ ^ _07_;
  assign _36_ = ~(_29_ ^ _11_);
  assign binary_o[6] = _36_ ^ _01_;
  assign _37_ = ~(_32_ ^ _13_);
  assign binary_o[7] = _37_ ^ _12_;
  assign binary_o[15] = gray_i[15];
  assign \scan_xor.i  = gray_i;
  assign \scan_xor.o  = { gray_i[15], binary_o[14:0] };
  assign \scan_xor.scanN.row[0].fill  = 16'h0000;
  assign \scan_xor.scanN.row[0].shifted  = { 1'h0, gray_i[15:1] };
  assign \scan_xor.scanN.row[1].fill  = 16'h0000;
  assign \scan_xor.scanN.row[1].shifted [15:12] = { 2'h0, gray_i[15], binary_o[14] };
  assign \scan_xor.scanN.row[2].fill  = 16'h0000;
  assign \scan_xor.scanN.row[2].shifted [15:8] = { 4'h0, gray_i[15], binary_o[14:12] };
  assign \scan_xor.scanN.row[3].fill  = 16'h0000;
  assign \scan_xor.scanN.row[3].shifted  = { 8'h00, gray_i[15], binary_o[14:8] };
  assign { \scan_xor.t [79:56], \scan_xor.t [47:36], \scan_xor.t [31:18], \scan_xor.t [15:0] } = { gray_i[15], binary_o[14:0], gray_i[15], binary_o[14:8], gray_i[15], binary_o[14:12], \scan_xor.scanN.row[2].shifted [7:0], gray_i[15], binary_o[14], \scan_xor.scanN.row[1].shifted [11:0], gray_i };
endmodule
