module bsg_mux_one_hot(data_i, sel_one_hot_i, data_o);
  input [15:0] data_i;
  wire [15:0] data_i;
  wire [15:0] data_masked;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire \reduce[0].gather ;
  wire \reduce[10].gather ;
  wire \reduce[11].gather ;
  wire \reduce[12].gather ;
  wire \reduce[13].gather ;
  wire \reduce[14].gather ;
  wire \reduce[15].gather ;
  wire \reduce[1].gather ;
  wire \reduce[2].gather ;
  wire \reduce[3].gather ;
  wire \reduce[4].gather ;
  wire \reduce[5].gather ;
  wire \reduce[6].gather ;
  wire \reduce[7].gather ;
  wire \reduce[8].gather ;
  wire \reduce[9].gather ;
  input sel_one_hot_i;
  wire sel_one_hot_i;
  assign \reduce[5].gather  = sel_one_hot_i & data_i[5];
  assign \reduce[6].gather  = data_i[6] & sel_one_hot_i;
  assign \reduce[7].gather  = data_i[7] & sel_one_hot_i;
  assign \reduce[8].gather  = data_i[8] & sel_one_hot_i;
  assign \reduce[9].gather  = data_i[9] & sel_one_hot_i;
  assign \reduce[10].gather  = data_i[10] & sel_one_hot_i;
  assign \reduce[11].gather  = data_i[11] & sel_one_hot_i;
  assign \reduce[12].gather  = data_i[12] & sel_one_hot_i;
  assign \reduce[13].gather  = data_i[13] & sel_one_hot_i;
  assign \reduce[14].gather  = data_i[14] & sel_one_hot_i;
  assign \reduce[15].gather  = data_i[15] & sel_one_hot_i;
  assign \reduce[0].gather  = data_i[0] & sel_one_hot_i;
  assign \reduce[1].gather  = data_i[1] & sel_one_hot_i;
  assign \reduce[2].gather  = data_i[2] & sel_one_hot_i;
  assign \reduce[3].gather  = data_i[3] & sel_one_hot_i;
  assign \reduce[4].gather  = data_i[4] & sel_one_hot_i;
  assign data_masked = { \reduce[15].gather , \reduce[14].gather , \reduce[13].gather , \reduce[12].gather , \reduce[11].gather , \reduce[10].gather , \reduce[9].gather , \reduce[8].gather , \reduce[7].gather , \reduce[6].gather , \reduce[5].gather , \reduce[4].gather , \reduce[3].gather , \reduce[2].gather , \reduce[1].gather , \reduce[0].gather  };
  assign data_o = { \reduce[15].gather , \reduce[14].gather , \reduce[13].gather , \reduce[12].gather , \reduce[11].gather , \reduce[10].gather , \reduce[9].gather , \reduce[8].gather , \reduce[7].gather , \reduce[6].gather , \reduce[5].gather , \reduce[4].gather , \reduce[3].gather , \reduce[2].gather , \reduce[1].gather , \reduce[0].gather  };
endmodule
