module bsg_crossbar_o_by_i(i, sel_oi_one_hot_i, o);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  input [255:0] i;
  wire [255:0] i;
  wire [255:0] \l[0].mux_one_hot.data_i ;
  wire [15:0] \l[0].mux_one_hot.data_o ;
  wire [15:0] \l[0].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[10].mux_one_hot.data_i ;
  wire [15:0] \l[10].mux_one_hot.data_o ;
  wire [15:0] \l[10].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[11].mux_one_hot.data_i ;
  wire [15:0] \l[11].mux_one_hot.data_o ;
  wire [15:0] \l[11].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[12].mux_one_hot.data_i ;
  wire [15:0] \l[12].mux_one_hot.data_o ;
  wire [15:0] \l[12].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[13].mux_one_hot.data_i ;
  wire [15:0] \l[13].mux_one_hot.data_o ;
  wire [15:0] \l[13].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[14].mux_one_hot.data_i ;
  wire [15:0] \l[14].mux_one_hot.data_o ;
  wire [15:0] \l[14].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[15].mux_one_hot.data_i ;
  wire [15:0] \l[15].mux_one_hot.data_o ;
  wire [15:0] \l[15].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[1].mux_one_hot.data_i ;
  wire [15:0] \l[1].mux_one_hot.data_o ;
  wire [15:0] \l[1].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[2].mux_one_hot.data_i ;
  wire [15:0] \l[2].mux_one_hot.data_o ;
  wire [15:0] \l[2].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[3].mux_one_hot.data_i ;
  wire [15:0] \l[3].mux_one_hot.data_o ;
  wire [15:0] \l[3].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[4].mux_one_hot.data_i ;
  wire [15:0] \l[4].mux_one_hot.data_o ;
  wire [15:0] \l[4].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[5].mux_one_hot.data_i ;
  wire [15:0] \l[5].mux_one_hot.data_o ;
  wire [15:0] \l[5].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[6].mux_one_hot.data_i ;
  wire [15:0] \l[6].mux_one_hot.data_o ;
  wire [15:0] \l[6].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[7].mux_one_hot.data_i ;
  wire [15:0] \l[7].mux_one_hot.data_o ;
  wire [15:0] \l[7].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[8].mux_one_hot.data_i ;
  wire [15:0] \l[8].mux_one_hot.data_o ;
  wire [15:0] \l[8].mux_one_hot.sel_one_hot_i ;
  wire [255:0] \l[9].mux_one_hot.data_i ;
  wire [15:0] \l[9].mux_one_hot.data_o ;
  wire [15:0] \l[9].mux_one_hot.sel_one_hot_i ;
  output [255:0] o;
  wire [255:0] o;
  input [255:0] sel_oi_one_hot_i;
  wire [255:0] sel_oi_one_hot_i;
  assign o[54] = _00675_ | _00660_;
  assign _00676_ = sel_oi_one_hot_i[48] & i[5];
  assign _00677_ = sel_oi_one_hot_i[49] & i[21];
  assign _00678_ = _00677_ | _00676_;
  assign _00679_ = sel_oi_one_hot_i[50] & i[37];
  assign _00680_ = sel_oi_one_hot_i[51] & i[53];
  assign _00681_ = _00680_ | _00679_;
  assign _00682_ = _00681_ | _00678_;
  assign _00683_ = sel_oi_one_hot_i[52] & i[69];
  assign _00684_ = sel_oi_one_hot_i[53] & i[85];
  assign _00685_ = _00684_ | _00683_;
  assign _00686_ = sel_oi_one_hot_i[54] & i[101];
  assign _00687_ = sel_oi_one_hot_i[55] & i[117];
  assign _00688_ = _00687_ | _00686_;
  assign _00689_ = _00688_ | _00685_;
  assign _00690_ = _00689_ | _00682_;
  assign _00691_ = sel_oi_one_hot_i[56] & i[133];
  assign _00692_ = sel_oi_one_hot_i[57] & i[149];
  assign _00693_ = _00692_ | _00691_;
  assign _00694_ = sel_oi_one_hot_i[58] & i[165];
  assign _00695_ = sel_oi_one_hot_i[59] & i[181];
  assign _00696_ = _00695_ | _00694_;
  assign _00697_ = _00696_ | _00693_;
  assign _00698_ = sel_oi_one_hot_i[60] & i[197];
  assign _00699_ = sel_oi_one_hot_i[61] & i[213];
  assign _00700_ = _00699_ | _00698_;
  assign _00701_ = sel_oi_one_hot_i[62] & i[229];
  assign _00702_ = sel_oi_one_hot_i[63] & i[245];
  assign _00703_ = _00702_ | _00701_;
  assign _00704_ = _00703_ | _00700_;
  assign _00705_ = _00704_ | _00697_;
  assign o[53] = _00705_ | _00690_;
  assign _00706_ = sel_oi_one_hot_i[48] & i[4];
  assign _00707_ = sel_oi_one_hot_i[49] & i[20];
  assign _00708_ = _00707_ | _00706_;
  assign _00709_ = sel_oi_one_hot_i[50] & i[36];
  assign _00710_ = sel_oi_one_hot_i[51] & i[52];
  assign _00711_ = _00710_ | _00709_;
  assign _00712_ = _00711_ | _00708_;
  assign _00713_ = sel_oi_one_hot_i[52] & i[68];
  assign _00714_ = sel_oi_one_hot_i[53] & i[84];
  assign _00715_ = _00714_ | _00713_;
  assign _00716_ = sel_oi_one_hot_i[54] & i[100];
  assign _00717_ = sel_oi_one_hot_i[55] & i[116];
  assign _00718_ = _00717_ | _00716_;
  assign _00719_ = _00718_ | _00715_;
  assign _00720_ = _00719_ | _00712_;
  assign _00721_ = sel_oi_one_hot_i[56] & i[132];
  assign _00722_ = sel_oi_one_hot_i[57] & i[148];
  assign _00723_ = _00722_ | _00721_;
  assign _00724_ = sel_oi_one_hot_i[58] & i[164];
  assign _00725_ = sel_oi_one_hot_i[59] & i[180];
  assign _00726_ = _00725_ | _00724_;
  assign _00727_ = _00726_ | _00723_;
  assign _00728_ = sel_oi_one_hot_i[60] & i[196];
  assign _00729_ = sel_oi_one_hot_i[61] & i[212];
  assign _00730_ = _00729_ | _00728_;
  assign _00731_ = sel_oi_one_hot_i[62] & i[228];
  assign _00732_ = sel_oi_one_hot_i[63] & i[244];
  assign _00733_ = _00732_ | _00731_;
  assign _00734_ = _00733_ | _00730_;
  assign _00735_ = _00734_ | _00727_;
  assign o[52] = _00735_ | _00720_;
  assign _00736_ = sel_oi_one_hot_i[48] & i[3];
  assign _00737_ = sel_oi_one_hot_i[49] & i[19];
  assign _00738_ = _00737_ | _00736_;
  assign _00739_ = sel_oi_one_hot_i[50] & i[35];
  assign _00740_ = sel_oi_one_hot_i[51] & i[51];
  assign _00741_ = _00740_ | _00739_;
  assign _00742_ = _00741_ | _00738_;
  assign _00743_ = sel_oi_one_hot_i[52] & i[67];
  assign _00744_ = sel_oi_one_hot_i[53] & i[83];
  assign _00745_ = _00744_ | _00743_;
  assign _00746_ = sel_oi_one_hot_i[54] & i[99];
  assign _00747_ = sel_oi_one_hot_i[55] & i[115];
  assign _00748_ = _00747_ | _00746_;
  assign _00749_ = _00748_ | _00745_;
  assign _00750_ = _00749_ | _00742_;
  assign _00751_ = sel_oi_one_hot_i[56] & i[131];
  assign _00752_ = sel_oi_one_hot_i[57] & i[147];
  assign _00753_ = _00752_ | _00751_;
  assign _00754_ = sel_oi_one_hot_i[58] & i[163];
  assign _00755_ = sel_oi_one_hot_i[59] & i[179];
  assign _00756_ = _00755_ | _00754_;
  assign _00757_ = _00756_ | _00753_;
  assign _00758_ = sel_oi_one_hot_i[60] & i[195];
  assign _00759_ = sel_oi_one_hot_i[61] & i[211];
  assign _00760_ = _00759_ | _00758_;
  assign _00761_ = sel_oi_one_hot_i[62] & i[227];
  assign _00762_ = sel_oi_one_hot_i[63] & i[243];
  assign _00763_ = _00762_ | _00761_;
  assign _00764_ = _00763_ | _00760_;
  assign _00765_ = _00764_ | _00757_;
  assign o[51] = _00765_ | _00750_;
  assign _00766_ = sel_oi_one_hot_i[0] & i[11];
  assign _00767_ = sel_oi_one_hot_i[1] & i[27];
  assign _00768_ = _00767_ | _00766_;
  assign _00769_ = sel_oi_one_hot_i[2] & i[43];
  assign _00770_ = sel_oi_one_hot_i[3] & i[59];
  assign _00771_ = _00770_ | _00769_;
  assign _00772_ = _00771_ | _00768_;
  assign _00773_ = sel_oi_one_hot_i[4] & i[75];
  assign _00774_ = sel_oi_one_hot_i[5] & i[91];
  assign _00775_ = _00774_ | _00773_;
  assign _00776_ = sel_oi_one_hot_i[6] & i[107];
  assign _00777_ = sel_oi_one_hot_i[7] & i[123];
  assign _00778_ = _00777_ | _00776_;
  assign _00779_ = _00778_ | _00775_;
  assign _00780_ = _00779_ | _00772_;
  assign _00781_ = sel_oi_one_hot_i[8] & i[139];
  assign _00782_ = sel_oi_one_hot_i[9] & i[155];
  assign _00783_ = _00782_ | _00781_;
  assign _00784_ = sel_oi_one_hot_i[10] & i[171];
  assign _00785_ = sel_oi_one_hot_i[11] & i[187];
  assign _00786_ = _00785_ | _00784_;
  assign _00787_ = _00786_ | _00783_;
  assign _00788_ = sel_oi_one_hot_i[12] & i[203];
  assign _00789_ = sel_oi_one_hot_i[13] & i[219];
  assign _00790_ = _00789_ | _00788_;
  assign _00791_ = sel_oi_one_hot_i[14] & i[235];
  assign _00792_ = sel_oi_one_hot_i[15] & i[251];
  assign _00793_ = _00792_ | _00791_;
  assign _00794_ = _00793_ | _00790_;
  assign _00795_ = _00794_ | _00787_;
  assign o[11] = _00795_ | _00780_;
  assign _00796_ = sel_oi_one_hot_i[48] & i[2];
  assign _00797_ = sel_oi_one_hot_i[49] & i[18];
  assign _00798_ = _00797_ | _00796_;
  assign _00799_ = sel_oi_one_hot_i[50] & i[34];
  assign _00800_ = sel_oi_one_hot_i[51] & i[50];
  assign _00801_ = _00800_ | _00799_;
  assign _00802_ = _00801_ | _00798_;
  assign _00803_ = sel_oi_one_hot_i[52] & i[66];
  assign _00804_ = sel_oi_one_hot_i[53] & i[82];
  assign _00805_ = _00804_ | _00803_;
  assign _00806_ = sel_oi_one_hot_i[54] & i[98];
  assign _00807_ = sel_oi_one_hot_i[55] & i[114];
  assign _00808_ = _00807_ | _00806_;
  assign _00809_ = _00808_ | _00805_;
  assign _00810_ = _00809_ | _00802_;
  assign _00811_ = sel_oi_one_hot_i[56] & i[130];
  assign _00812_ = sel_oi_one_hot_i[57] & i[146];
  assign _00813_ = _00812_ | _00811_;
  assign _00814_ = sel_oi_one_hot_i[58] & i[162];
  assign _00815_ = sel_oi_one_hot_i[59] & i[178];
  assign _00816_ = _00815_ | _00814_;
  assign _00817_ = _00816_ | _00813_;
  assign _00818_ = sel_oi_one_hot_i[60] & i[194];
  assign _00819_ = sel_oi_one_hot_i[61] & i[210];
  assign _00820_ = _00819_ | _00818_;
  assign _00821_ = sel_oi_one_hot_i[62] & i[226];
  assign _00822_ = sel_oi_one_hot_i[63] & i[242];
  assign _00823_ = _00822_ | _00821_;
  assign _00824_ = _00823_ | _00820_;
  assign _00825_ = _00824_ | _00817_;
  assign o[50] = _00825_ | _00810_;
  assign _00826_ = sel_oi_one_hot_i[48] & i[1];
  assign _00827_ = sel_oi_one_hot_i[49] & i[17];
  assign _00828_ = _00827_ | _00826_;
  assign _00829_ = sel_oi_one_hot_i[50] & i[33];
  assign _00830_ = sel_oi_one_hot_i[51] & i[49];
  assign _00831_ = _00830_ | _00829_;
  assign _00832_ = _00831_ | _00828_;
  assign _00833_ = sel_oi_one_hot_i[52] & i[65];
  assign _00834_ = sel_oi_one_hot_i[53] & i[81];
  assign _00835_ = _00834_ | _00833_;
  assign _00836_ = sel_oi_one_hot_i[54] & i[97];
  assign _00837_ = sel_oi_one_hot_i[55] & i[113];
  assign _00838_ = _00837_ | _00836_;
  assign _00839_ = _00838_ | _00835_;
  assign _00840_ = _00839_ | _00832_;
  assign _00841_ = sel_oi_one_hot_i[56] & i[129];
  assign _00842_ = sel_oi_one_hot_i[57] & i[145];
  assign _00843_ = _00842_ | _00841_;
  assign _00844_ = sel_oi_one_hot_i[58] & i[161];
  assign _00845_ = sel_oi_one_hot_i[59] & i[177];
  assign _00846_ = _00845_ | _00844_;
  assign _00847_ = _00846_ | _00843_;
  assign _00848_ = sel_oi_one_hot_i[60] & i[193];
  assign _00849_ = sel_oi_one_hot_i[61] & i[209];
  assign _00850_ = _00849_ | _00848_;
  assign _00851_ = sel_oi_one_hot_i[62] & i[225];
  assign _00852_ = sel_oi_one_hot_i[63] & i[241];
  assign _00853_ = _00852_ | _00851_;
  assign _00854_ = _00853_ | _00850_;
  assign _00855_ = _00854_ | _00847_;
  assign o[49] = _00855_ | _00840_;
  assign _00856_ = sel_oi_one_hot_i[48] & i[0];
  assign _00857_ = sel_oi_one_hot_i[49] & i[16];
  assign _00858_ = _00857_ | _00856_;
  assign _00859_ = sel_oi_one_hot_i[50] & i[32];
  assign _00860_ = sel_oi_one_hot_i[51] & i[48];
  assign _00861_ = _00860_ | _00859_;
  assign _00862_ = _00861_ | _00858_;
  assign _00863_ = sel_oi_one_hot_i[52] & i[64];
  assign _00864_ = sel_oi_one_hot_i[53] & i[80];
  assign _00865_ = _00864_ | _00863_;
  assign _00866_ = sel_oi_one_hot_i[54] & i[96];
  assign _00867_ = sel_oi_one_hot_i[55] & i[112];
  assign _00868_ = _00867_ | _00866_;
  assign _00869_ = _00868_ | _00865_;
  assign _00870_ = _00869_ | _00862_;
  assign _00871_ = sel_oi_one_hot_i[56] & i[128];
  assign _00872_ = sel_oi_one_hot_i[57] & i[144];
  assign _00873_ = _00872_ | _00871_;
  assign _00874_ = sel_oi_one_hot_i[58] & i[160];
  assign _00875_ = sel_oi_one_hot_i[59] & i[176];
  assign _00876_ = _00875_ | _00874_;
  assign _00877_ = _00876_ | _00873_;
  assign _00878_ = sel_oi_one_hot_i[60] & i[192];
  assign _00879_ = sel_oi_one_hot_i[61] & i[208];
  assign _00880_ = _00879_ | _00878_;
  assign _00881_ = sel_oi_one_hot_i[62] & i[224];
  assign _00882_ = sel_oi_one_hot_i[63] & i[240];
  assign _00883_ = _00882_ | _00881_;
  assign _00884_ = _00883_ | _00880_;
  assign _00885_ = _00884_ | _00877_;
  assign o[48] = _00885_ | _00870_;
  assign _00886_ = sel_oi_one_hot_i[0] & i[10];
  assign _00887_ = sel_oi_one_hot_i[1] & i[26];
  assign _00888_ = _00887_ | _00886_;
  assign _00889_ = sel_oi_one_hot_i[2] & i[42];
  assign _00890_ = sel_oi_one_hot_i[3] & i[58];
  assign _00891_ = _00890_ | _00889_;
  assign _00892_ = _00891_ | _00888_;
  assign _00893_ = sel_oi_one_hot_i[4] & i[74];
  assign _00894_ = sel_oi_one_hot_i[5] & i[90];
  assign _00895_ = _00894_ | _00893_;
  assign _00896_ = sel_oi_one_hot_i[6] & i[106];
  assign _00897_ = sel_oi_one_hot_i[7] & i[122];
  assign _00898_ = _00897_ | _00896_;
  assign _00899_ = _00898_ | _00895_;
  assign _00900_ = _00899_ | _00892_;
  assign _00901_ = sel_oi_one_hot_i[8] & i[138];
  assign _00902_ = sel_oi_one_hot_i[9] & i[154];
  assign _00903_ = _00902_ | _00901_;
  assign _00904_ = sel_oi_one_hot_i[10] & i[170];
  assign _00905_ = sel_oi_one_hot_i[11] & i[186];
  assign _00906_ = _00905_ | _00904_;
  assign _00907_ = _00906_ | _00903_;
  assign _00908_ = sel_oi_one_hot_i[12] & i[202];
  assign _00909_ = sel_oi_one_hot_i[13] & i[218];
  assign _00910_ = _00909_ | _00908_;
  assign _00911_ = sel_oi_one_hot_i[14] & i[234];
  assign _00912_ = sel_oi_one_hot_i[15] & i[250];
  assign _00913_ = _00912_ | _00911_;
  assign _00914_ = _00913_ | _00910_;
  assign _00915_ = _00914_ | _00907_;
  assign o[10] = _00915_ | _00900_;
  assign _00916_ = sel_oi_one_hot_i[64] & i[15];
  assign _00917_ = sel_oi_one_hot_i[65] & i[31];
  assign _00918_ = _00917_ | _00916_;
  assign _00919_ = sel_oi_one_hot_i[66] & i[47];
  assign _00920_ = sel_oi_one_hot_i[67] & i[63];
  assign _00921_ = _00920_ | _00919_;
  assign _00922_ = _00921_ | _00918_;
  assign _00923_ = sel_oi_one_hot_i[68] & i[79];
  assign _00924_ = sel_oi_one_hot_i[69] & i[95];
  assign _00925_ = _00924_ | _00923_;
  assign _00926_ = sel_oi_one_hot_i[70] & i[111];
  assign _00927_ = sel_oi_one_hot_i[71] & i[127];
  assign _00928_ = _00927_ | _00926_;
  assign _00929_ = _00928_ | _00925_;
  assign _00930_ = _00929_ | _00922_;
  assign _00931_ = sel_oi_one_hot_i[72] & i[143];
  assign _00932_ = sel_oi_one_hot_i[73] & i[159];
  assign _00933_ = _00932_ | _00931_;
  assign _00934_ = sel_oi_one_hot_i[74] & i[175];
  assign _00935_ = sel_oi_one_hot_i[75] & i[191];
  assign _00936_ = _00935_ | _00934_;
  assign _00937_ = _00936_ | _00933_;
  assign _00938_ = sel_oi_one_hot_i[76] & i[207];
  assign _00939_ = sel_oi_one_hot_i[77] & i[223];
  assign _00940_ = _00939_ | _00938_;
  assign _00941_ = sel_oi_one_hot_i[78] & i[239];
  assign _00942_ = sel_oi_one_hot_i[79] & i[255];
  assign _00943_ = _00942_ | _00941_;
  assign _00944_ = _00943_ | _00940_;
  assign _00945_ = _00944_ | _00937_;
  assign o[79] = _00945_ | _00930_;
  assign _00946_ = sel_oi_one_hot_i[64] & i[14];
  assign _00947_ = sel_oi_one_hot_i[65] & i[30];
  assign _00948_ = _00947_ | _00946_;
  assign _00949_ = sel_oi_one_hot_i[66] & i[46];
  assign _00950_ = sel_oi_one_hot_i[67] & i[62];
  assign _00951_ = _00950_ | _00949_;
  assign _00952_ = _00951_ | _00948_;
  assign _00953_ = sel_oi_one_hot_i[68] & i[78];
  assign _00954_ = sel_oi_one_hot_i[69] & i[94];
  assign _00955_ = _00954_ | _00953_;
  assign _00956_ = sel_oi_one_hot_i[70] & i[110];
  assign _00957_ = sel_oi_one_hot_i[71] & i[126];
  assign _00958_ = _00957_ | _00956_;
  assign _00959_ = _00958_ | _00955_;
  assign _00960_ = _00959_ | _00952_;
  assign _00961_ = sel_oi_one_hot_i[72] & i[142];
  assign _00962_ = sel_oi_one_hot_i[73] & i[158];
  assign _00963_ = _00962_ | _00961_;
  assign _00964_ = sel_oi_one_hot_i[74] & i[174];
  assign _00965_ = sel_oi_one_hot_i[75] & i[190];
  assign _00966_ = _00965_ | _00964_;
  assign _00967_ = _00966_ | _00963_;
  assign _00968_ = sel_oi_one_hot_i[76] & i[206];
  assign _00969_ = sel_oi_one_hot_i[77] & i[222];
  assign _00970_ = _00969_ | _00968_;
  assign _00971_ = sel_oi_one_hot_i[78] & i[238];
  assign _00972_ = sel_oi_one_hot_i[79] & i[254];
  assign _00973_ = _00972_ | _00971_;
  assign _00974_ = _00973_ | _00970_;
  assign _00975_ = _00974_ | _00967_;
  assign o[78] = _00975_ | _00960_;
  assign _00976_ = sel_oi_one_hot_i[64] & i[13];
  assign _00977_ = sel_oi_one_hot_i[65] & i[29];
  assign _00978_ = _00977_ | _00976_;
  assign _00979_ = sel_oi_one_hot_i[66] & i[45];
  assign _00980_ = sel_oi_one_hot_i[67] & i[61];
  assign _00981_ = _00980_ | _00979_;
  assign _00982_ = _00981_ | _00978_;
  assign _00983_ = sel_oi_one_hot_i[68] & i[77];
  assign _00984_ = sel_oi_one_hot_i[69] & i[93];
  assign _00985_ = _00984_ | _00983_;
  assign _00986_ = sel_oi_one_hot_i[70] & i[109];
  assign _00987_ = sel_oi_one_hot_i[71] & i[125];
  assign _00988_ = _00987_ | _00986_;
  assign _00989_ = _00988_ | _00985_;
  assign _00990_ = _00989_ | _00982_;
  assign _00991_ = sel_oi_one_hot_i[72] & i[141];
  assign _00992_ = sel_oi_one_hot_i[73] & i[157];
  assign _00993_ = _00992_ | _00991_;
  assign _00994_ = sel_oi_one_hot_i[74] & i[173];
  assign _00995_ = sel_oi_one_hot_i[75] & i[189];
  assign _00996_ = _00995_ | _00994_;
  assign _00997_ = _00996_ | _00993_;
  assign _00998_ = sel_oi_one_hot_i[76] & i[205];
  assign _00999_ = sel_oi_one_hot_i[77] & i[221];
  assign _01000_ = _00999_ | _00998_;
  assign _01001_ = sel_oi_one_hot_i[78] & i[237];
  assign _01002_ = sel_oi_one_hot_i[79] & i[253];
  assign _01003_ = _01002_ | _01001_;
  assign _01004_ = _01003_ | _01000_;
  assign _01005_ = _01004_ | _00997_;
  assign o[77] = _01005_ | _00990_;
  assign _01006_ = sel_oi_one_hot_i[0] & i[9];
  assign _01007_ = sel_oi_one_hot_i[1] & i[25];
  assign _01008_ = _01007_ | _01006_;
  assign _01009_ = sel_oi_one_hot_i[2] & i[41];
  assign _01010_ = sel_oi_one_hot_i[3] & i[57];
  assign _01011_ = _01010_ | _01009_;
  assign _01012_ = _01011_ | _01008_;
  assign _01013_ = sel_oi_one_hot_i[4] & i[73];
  assign _01014_ = sel_oi_one_hot_i[5] & i[89];
  assign _01015_ = _01014_ | _01013_;
  assign _01016_ = sel_oi_one_hot_i[6] & i[105];
  assign _01017_ = sel_oi_one_hot_i[7] & i[121];
  assign _01018_ = _01017_ | _01016_;
  assign _01019_ = _01018_ | _01015_;
  assign _01020_ = _01019_ | _01012_;
  assign _01021_ = sel_oi_one_hot_i[8] & i[137];
  assign _01022_ = sel_oi_one_hot_i[9] & i[153];
  assign _01023_ = _01022_ | _01021_;
  assign _01024_ = sel_oi_one_hot_i[10] & i[169];
  assign _01025_ = sel_oi_one_hot_i[11] & i[185];
  assign _01026_ = _01025_ | _01024_;
  assign _01027_ = _01026_ | _01023_;
  assign _01028_ = sel_oi_one_hot_i[12] & i[201];
  assign _01029_ = sel_oi_one_hot_i[13] & i[217];
  assign _01030_ = _01029_ | _01028_;
  assign _01031_ = sel_oi_one_hot_i[14] & i[233];
  assign _01032_ = sel_oi_one_hot_i[15] & i[249];
  assign _01033_ = _01032_ | _01031_;
  assign _01034_ = _01033_ | _01030_;
  assign _01035_ = _01034_ | _01027_;
  assign o[9] = _01035_ | _01020_;
  assign _01036_ = sel_oi_one_hot_i[64] & i[12];
  assign _01037_ = sel_oi_one_hot_i[65] & i[28];
  assign _01038_ = _01037_ | _01036_;
  assign _01039_ = sel_oi_one_hot_i[66] & i[44];
  assign _01040_ = sel_oi_one_hot_i[67] & i[60];
  assign _01041_ = _01040_ | _01039_;
  assign _01042_ = _01041_ | _01038_;
  assign _01043_ = sel_oi_one_hot_i[68] & i[76];
  assign _01044_ = sel_oi_one_hot_i[69] & i[92];
  assign _01045_ = _01044_ | _01043_;
  assign _01046_ = sel_oi_one_hot_i[70] & i[108];
  assign _01047_ = sel_oi_one_hot_i[71] & i[124];
  assign _01048_ = _01047_ | _01046_;
  assign _01049_ = _01048_ | _01045_;
  assign _01050_ = _01049_ | _01042_;
  assign _01051_ = sel_oi_one_hot_i[72] & i[140];
  assign _01052_ = sel_oi_one_hot_i[73] & i[156];
  assign _01053_ = _01052_ | _01051_;
  assign _01054_ = sel_oi_one_hot_i[74] & i[172];
  assign _01055_ = sel_oi_one_hot_i[75] & i[188];
  assign _01056_ = _01055_ | _01054_;
  assign _01057_ = _01056_ | _01053_;
  assign _01058_ = sel_oi_one_hot_i[76] & i[204];
  assign _01059_ = sel_oi_one_hot_i[77] & i[220];
  assign _01060_ = _01059_ | _01058_;
  assign _01061_ = sel_oi_one_hot_i[78] & i[236];
  assign _01062_ = sel_oi_one_hot_i[79] & i[252];
  assign _01063_ = _01062_ | _01061_;
  assign _01064_ = _01063_ | _01060_;
  assign _01065_ = _01064_ | _01057_;
  assign o[76] = _01065_ | _01050_;
  assign _01066_ = sel_oi_one_hot_i[64] & i[11];
  assign _01067_ = sel_oi_one_hot_i[65] & i[27];
  assign _01068_ = _01067_ | _01066_;
  assign _01069_ = sel_oi_one_hot_i[66] & i[43];
  assign _01070_ = sel_oi_one_hot_i[67] & i[59];
  assign _01071_ = _01070_ | _01069_;
  assign _01072_ = _01071_ | _01068_;
  assign _01073_ = sel_oi_one_hot_i[68] & i[75];
  assign _01074_ = sel_oi_one_hot_i[69] & i[91];
  assign _01075_ = _01074_ | _01073_;
  assign _01076_ = sel_oi_one_hot_i[70] & i[107];
  assign _01077_ = sel_oi_one_hot_i[71] & i[123];
  assign _01078_ = _01077_ | _01076_;
  assign _01079_ = _01078_ | _01075_;
  assign _01080_ = _01079_ | _01072_;
  assign _01081_ = sel_oi_one_hot_i[72] & i[139];
  assign _01082_ = sel_oi_one_hot_i[73] & i[155];
  assign _01083_ = _01082_ | _01081_;
  assign _01084_ = sel_oi_one_hot_i[74] & i[171];
  assign _01085_ = sel_oi_one_hot_i[75] & i[187];
  assign _01086_ = _01085_ | _01084_;
  assign _01087_ = _01086_ | _01083_;
  assign _01088_ = sel_oi_one_hot_i[76] & i[203];
  assign _01089_ = sel_oi_one_hot_i[77] & i[219];
  assign _01090_ = _01089_ | _01088_;
  assign _01091_ = sel_oi_one_hot_i[78] & i[235];
  assign _01092_ = sel_oi_one_hot_i[79] & i[251];
  assign _01093_ = _01092_ | _01091_;
  assign _01094_ = _01093_ | _01090_;
  assign _01095_ = _01094_ | _01087_;
  assign o[75] = _01095_ | _01080_;
  assign _01096_ = sel_oi_one_hot_i[64] & i[10];
  assign _01097_ = sel_oi_one_hot_i[65] & i[26];
  assign _01098_ = _01097_ | _01096_;
  assign _01099_ = sel_oi_one_hot_i[66] & i[42];
  assign _01100_ = sel_oi_one_hot_i[67] & i[58];
  assign _01101_ = _01100_ | _01099_;
  assign _01102_ = _01101_ | _01098_;
  assign _01103_ = sel_oi_one_hot_i[68] & i[74];
  assign _01104_ = sel_oi_one_hot_i[69] & i[90];
  assign _01105_ = _01104_ | _01103_;
  assign _01106_ = sel_oi_one_hot_i[70] & i[106];
  assign _01107_ = sel_oi_one_hot_i[71] & i[122];
  assign _01108_ = _01107_ | _01106_;
  assign _01109_ = _01108_ | _01105_;
  assign _01110_ = _01109_ | _01102_;
  assign _01111_ = sel_oi_one_hot_i[72] & i[138];
  assign _01112_ = sel_oi_one_hot_i[73] & i[154];
  assign _01113_ = _01112_ | _01111_;
  assign _01114_ = sel_oi_one_hot_i[74] & i[170];
  assign _01115_ = sel_oi_one_hot_i[75] & i[186];
  assign _01116_ = _01115_ | _01114_;
  assign _01117_ = _01116_ | _01113_;
  assign _01118_ = sel_oi_one_hot_i[76] & i[202];
  assign _01119_ = sel_oi_one_hot_i[77] & i[218];
  assign _01120_ = _01119_ | _01118_;
  assign _01121_ = sel_oi_one_hot_i[78] & i[234];
  assign _01122_ = sel_oi_one_hot_i[79] & i[250];
  assign _01123_ = _01122_ | _01121_;
  assign _01124_ = _01123_ | _01120_;
  assign _01125_ = _01124_ | _01117_;
  assign o[74] = _01125_ | _01110_;
  assign _01126_ = sel_oi_one_hot_i[64] & i[9];
  assign _01127_ = sel_oi_one_hot_i[65] & i[25];
  assign _01128_ = _01127_ | _01126_;
  assign _01129_ = sel_oi_one_hot_i[66] & i[41];
  assign _01130_ = sel_oi_one_hot_i[67] & i[57];
  assign _01131_ = _01130_ | _01129_;
  assign _01132_ = _01131_ | _01128_;
  assign _01133_ = sel_oi_one_hot_i[68] & i[73];
  assign _01134_ = sel_oi_one_hot_i[69] & i[89];
  assign _01135_ = _01134_ | _01133_;
  assign _01136_ = sel_oi_one_hot_i[70] & i[105];
  assign _01137_ = sel_oi_one_hot_i[71] & i[121];
  assign _01138_ = _01137_ | _01136_;
  assign _01139_ = _01138_ | _01135_;
  assign _01140_ = _01139_ | _01132_;
  assign _01141_ = sel_oi_one_hot_i[72] & i[137];
  assign _01142_ = sel_oi_one_hot_i[73] & i[153];
  assign _01143_ = _01142_ | _01141_;
  assign _01144_ = sel_oi_one_hot_i[74] & i[169];
  assign _01145_ = sel_oi_one_hot_i[75] & i[185];
  assign _01146_ = _01145_ | _01144_;
  assign _01147_ = _01146_ | _01143_;
  assign _01148_ = sel_oi_one_hot_i[76] & i[201];
  assign _01149_ = sel_oi_one_hot_i[77] & i[217];
  assign _01150_ = _01149_ | _01148_;
  assign _01151_ = sel_oi_one_hot_i[78] & i[233];
  assign _01152_ = sel_oi_one_hot_i[79] & i[249];
  assign _01153_ = _01152_ | _01151_;
  assign _01154_ = _01153_ | _01150_;
  assign _01155_ = _01154_ | _01147_;
  assign o[73] = _01155_ | _01140_;
  assign _01156_ = sel_oi_one_hot_i[64] & i[8];
  assign _01157_ = sel_oi_one_hot_i[65] & i[24];
  assign _01158_ = _01157_ | _01156_;
  assign _01159_ = sel_oi_one_hot_i[66] & i[40];
  assign _01160_ = sel_oi_one_hot_i[67] & i[56];
  assign _01161_ = _01160_ | _01159_;
  assign _01162_ = _01161_ | _01158_;
  assign _01163_ = sel_oi_one_hot_i[68] & i[72];
  assign _01164_ = sel_oi_one_hot_i[69] & i[88];
  assign _01165_ = _01164_ | _01163_;
  assign _01166_ = sel_oi_one_hot_i[70] & i[104];
  assign _01167_ = sel_oi_one_hot_i[71] & i[120];
  assign _01168_ = _01167_ | _01166_;
  assign _01169_ = _01168_ | _01165_;
  assign _01170_ = _01169_ | _01162_;
  assign _01171_ = sel_oi_one_hot_i[72] & i[136];
  assign _01172_ = sel_oi_one_hot_i[73] & i[152];
  assign _01173_ = _01172_ | _01171_;
  assign _01174_ = sel_oi_one_hot_i[74] & i[168];
  assign _01175_ = sel_oi_one_hot_i[75] & i[184];
  assign _01176_ = _01175_ | _01174_;
  assign _01177_ = _01176_ | _01173_;
  assign _01178_ = sel_oi_one_hot_i[76] & i[200];
  assign _01179_ = sel_oi_one_hot_i[77] & i[216];
  assign _01180_ = _01179_ | _01178_;
  assign _01181_ = sel_oi_one_hot_i[78] & i[232];
  assign _01182_ = sel_oi_one_hot_i[79] & i[248];
  assign _01183_ = _01182_ | _01181_;
  assign _01184_ = _01183_ | _01180_;
  assign _01185_ = _01184_ | _01177_;
  assign o[72] = _01185_ | _01170_;
  assign _01186_ = sel_oi_one_hot_i[64] & i[7];
  assign _01187_ = sel_oi_one_hot_i[65] & i[23];
  assign _01188_ = _01187_ | _01186_;
  assign _01189_ = sel_oi_one_hot_i[66] & i[39];
  assign _01190_ = sel_oi_one_hot_i[67] & i[55];
  assign _01191_ = _01190_ | _01189_;
  assign _01192_ = _01191_ | _01188_;
  assign _01193_ = sel_oi_one_hot_i[68] & i[71];
  assign _01194_ = sel_oi_one_hot_i[69] & i[87];
  assign _01195_ = _01194_ | _01193_;
  assign _01196_ = sel_oi_one_hot_i[70] & i[103];
  assign _01197_ = sel_oi_one_hot_i[71] & i[119];
  assign _01198_ = _01197_ | _01196_;
  assign _01199_ = _01198_ | _01195_;
  assign _01200_ = _01199_ | _01192_;
  assign _01201_ = sel_oi_one_hot_i[72] & i[135];
  assign _01202_ = sel_oi_one_hot_i[73] & i[151];
  assign _01203_ = _01202_ | _01201_;
  assign _01204_ = sel_oi_one_hot_i[74] & i[167];
  assign _01205_ = sel_oi_one_hot_i[75] & i[183];
  assign _01206_ = _01205_ | _01204_;
  assign _01207_ = _01206_ | _01203_;
  assign _01208_ = sel_oi_one_hot_i[76] & i[199];
  assign _01209_ = sel_oi_one_hot_i[77] & i[215];
  assign _01210_ = _01209_ | _01208_;
  assign _01211_ = sel_oi_one_hot_i[78] & i[231];
  assign _01212_ = sel_oi_one_hot_i[79] & i[247];
  assign _01213_ = _01212_ | _01211_;
  assign _01214_ = _01213_ | _01210_;
  assign _01215_ = _01214_ | _01207_;
  assign o[71] = _01215_ | _01200_;
  assign _01216_ = sel_oi_one_hot_i[64] & i[6];
  assign _01217_ = sel_oi_one_hot_i[65] & i[22];
  assign _01218_ = _01217_ | _01216_;
  assign _01219_ = sel_oi_one_hot_i[66] & i[38];
  assign _01220_ = sel_oi_one_hot_i[67] & i[54];
  assign _01221_ = _01220_ | _01219_;
  assign _01222_ = _01221_ | _01218_;
  assign _01223_ = sel_oi_one_hot_i[68] & i[70];
  assign _01224_ = sel_oi_one_hot_i[69] & i[86];
  assign _01225_ = _01224_ | _01223_;
  assign _01226_ = sel_oi_one_hot_i[70] & i[102];
  assign _01227_ = sel_oi_one_hot_i[71] & i[118];
  assign _01228_ = _01227_ | _01226_;
  assign _01229_ = _01228_ | _01225_;
  assign _01230_ = _01229_ | _01222_;
  assign _01231_ = sel_oi_one_hot_i[72] & i[134];
  assign _01232_ = sel_oi_one_hot_i[73] & i[150];
  assign _01233_ = _01232_ | _01231_;
  assign _01234_ = sel_oi_one_hot_i[74] & i[166];
  assign _01235_ = sel_oi_one_hot_i[75] & i[182];
  assign _01236_ = _01235_ | _01234_;
  assign _01237_ = _01236_ | _01233_;
  assign _01238_ = sel_oi_one_hot_i[76] & i[198];
  assign _01239_ = sel_oi_one_hot_i[77] & i[214];
  assign _01240_ = _01239_ | _01238_;
  assign _01241_ = sel_oi_one_hot_i[78] & i[230];
  assign _01242_ = sel_oi_one_hot_i[79] & i[246];
  assign _01243_ = _01242_ | _01241_;
  assign _01244_ = _01243_ | _01240_;
  assign _01245_ = _01244_ | _01237_;
  assign o[70] = _01245_ | _01230_;
  assign _01246_ = sel_oi_one_hot_i[64] & i[5];
  assign _01247_ = sel_oi_one_hot_i[65] & i[21];
  assign _01248_ = _01247_ | _01246_;
  assign _01249_ = sel_oi_one_hot_i[66] & i[37];
  assign _01250_ = sel_oi_one_hot_i[67] & i[53];
  assign _01251_ = _01250_ | _01249_;
  assign _01252_ = _01251_ | _01248_;
  assign _01253_ = sel_oi_one_hot_i[68] & i[69];
  assign _01254_ = sel_oi_one_hot_i[69] & i[85];
  assign _01255_ = _01254_ | _01253_;
  assign _01256_ = sel_oi_one_hot_i[70] & i[101];
  assign _01257_ = sel_oi_one_hot_i[71] & i[117];
  assign _01258_ = _01257_ | _01256_;
  assign _01259_ = _01258_ | _01255_;
  assign _01260_ = _01259_ | _01252_;
  assign _01261_ = sel_oi_one_hot_i[72] & i[133];
  assign _01262_ = sel_oi_one_hot_i[73] & i[149];
  assign _01263_ = _01262_ | _01261_;
  assign _01264_ = sel_oi_one_hot_i[74] & i[165];
  assign _01265_ = sel_oi_one_hot_i[75] & i[181];
  assign _01266_ = _01265_ | _01264_;
  assign _01267_ = _01266_ | _01263_;
  assign _01268_ = sel_oi_one_hot_i[76] & i[197];
  assign _01269_ = sel_oi_one_hot_i[77] & i[213];
  assign _01270_ = _01269_ | _01268_;
  assign _01271_ = sel_oi_one_hot_i[78] & i[229];
  assign _01272_ = sel_oi_one_hot_i[79] & i[245];
  assign _01273_ = _01272_ | _01271_;
  assign _01274_ = _01273_ | _01270_;
  assign _01275_ = _01274_ | _01267_;
  assign o[69] = _01275_ | _01260_;
  assign _01276_ = sel_oi_one_hot_i[64] & i[4];
  assign _01277_ = sel_oi_one_hot_i[65] & i[20];
  assign _01278_ = _01277_ | _01276_;
  assign _01279_ = sel_oi_one_hot_i[66] & i[36];
  assign _01280_ = sel_oi_one_hot_i[67] & i[52];
  assign _01281_ = _01280_ | _01279_;
  assign _01282_ = _01281_ | _01278_;
  assign _01283_ = sel_oi_one_hot_i[68] & i[68];
  assign _01284_ = sel_oi_one_hot_i[69] & i[84];
  assign _01285_ = _01284_ | _01283_;
  assign _01286_ = sel_oi_one_hot_i[70] & i[100];
  assign _01287_ = sel_oi_one_hot_i[71] & i[116];
  assign _01288_ = _01287_ | _01286_;
  assign _01289_ = _01288_ | _01285_;
  assign _01290_ = _01289_ | _01282_;
  assign _01291_ = sel_oi_one_hot_i[72] & i[132];
  assign _01292_ = sel_oi_one_hot_i[73] & i[148];
  assign _01293_ = _01292_ | _01291_;
  assign _01294_ = sel_oi_one_hot_i[74] & i[164];
  assign _01295_ = sel_oi_one_hot_i[75] & i[180];
  assign _01296_ = _01295_ | _01294_;
  assign _01297_ = _01296_ | _01293_;
  assign _01298_ = sel_oi_one_hot_i[76] & i[196];
  assign _01299_ = sel_oi_one_hot_i[77] & i[212];
  assign _01300_ = _01299_ | _01298_;
  assign _01301_ = sel_oi_one_hot_i[78] & i[228];
  assign _01302_ = sel_oi_one_hot_i[79] & i[244];
  assign _01303_ = _01302_ | _01301_;
  assign _01304_ = _01303_ | _01300_;
  assign _01305_ = _01304_ | _01297_;
  assign o[68] = _01305_ | _01290_;
  assign _01306_ = sel_oi_one_hot_i[64] & i[3];
  assign _01307_ = sel_oi_one_hot_i[65] & i[19];
  assign _01308_ = _01307_ | _01306_;
  assign _01309_ = sel_oi_one_hot_i[66] & i[35];
  assign _01310_ = sel_oi_one_hot_i[67] & i[51];
  assign _01311_ = _01310_ | _01309_;
  assign _01312_ = _01311_ | _01308_;
  assign _01313_ = sel_oi_one_hot_i[68] & i[67];
  assign _01314_ = sel_oi_one_hot_i[69] & i[83];
  assign _01315_ = _01314_ | _01313_;
  assign _01316_ = sel_oi_one_hot_i[70] & i[99];
  assign _01317_ = sel_oi_one_hot_i[71] & i[115];
  assign _01318_ = _01317_ | _01316_;
  assign _01319_ = _01318_ | _01315_;
  assign _01320_ = _01319_ | _01312_;
  assign _01321_ = sel_oi_one_hot_i[72] & i[131];
  assign _01322_ = sel_oi_one_hot_i[73] & i[147];
  assign _01323_ = _01322_ | _01321_;
  assign _01324_ = sel_oi_one_hot_i[74] & i[163];
  assign _01325_ = sel_oi_one_hot_i[75] & i[179];
  assign _01326_ = _01325_ | _01324_;
  assign _01327_ = _01326_ | _01323_;
  assign _01328_ = sel_oi_one_hot_i[76] & i[195];
  assign _01329_ = sel_oi_one_hot_i[77] & i[211];
  assign _01330_ = _01329_ | _01328_;
  assign _01331_ = sel_oi_one_hot_i[78] & i[227];
  assign _01332_ = sel_oi_one_hot_i[79] & i[243];
  assign _01333_ = _01332_ | _01331_;
  assign _01334_ = _01333_ | _01330_;
  assign _01335_ = _01334_ | _01327_;
  assign o[67] = _01335_ | _01320_;
  assign _01336_ = sel_oi_one_hot_i[0] & i[8];
  assign _01337_ = sel_oi_one_hot_i[1] & i[24];
  assign _01338_ = _01337_ | _01336_;
  assign _01339_ = sel_oi_one_hot_i[2] & i[40];
  assign _01340_ = sel_oi_one_hot_i[3] & i[56];
  assign _01341_ = _01340_ | _01339_;
  assign _01342_ = _01341_ | _01338_;
  assign _01343_ = sel_oi_one_hot_i[4] & i[72];
  assign _01344_ = sel_oi_one_hot_i[5] & i[88];
  assign _01345_ = _01344_ | _01343_;
  assign _01346_ = sel_oi_one_hot_i[6] & i[104];
  assign _01347_ = sel_oi_one_hot_i[7] & i[120];
  assign _01348_ = _01347_ | _01346_;
  assign _01349_ = _01348_ | _01345_;
  assign _01350_ = _01349_ | _01342_;
  assign _01351_ = sel_oi_one_hot_i[8] & i[136];
  assign _01352_ = sel_oi_one_hot_i[9] & i[152];
  assign _01353_ = _01352_ | _01351_;
  assign _01354_ = sel_oi_one_hot_i[10] & i[168];
  assign _01355_ = sel_oi_one_hot_i[11] & i[184];
  assign _01356_ = _01355_ | _01354_;
  assign _01357_ = _01356_ | _01353_;
  assign _01358_ = sel_oi_one_hot_i[12] & i[200];
  assign _01359_ = sel_oi_one_hot_i[13] & i[216];
  assign _01360_ = _01359_ | _01358_;
  assign _01361_ = sel_oi_one_hot_i[14] & i[232];
  assign _01362_ = sel_oi_one_hot_i[15] & i[248];
  assign _01363_ = _01362_ | _01361_;
  assign _01364_ = _01363_ | _01360_;
  assign _01365_ = _01364_ | _01357_;
  assign o[8] = _01365_ | _01350_;
  assign _01366_ = sel_oi_one_hot_i[64] & i[2];
  assign _01367_ = sel_oi_one_hot_i[65] & i[18];
  assign _01368_ = _01367_ | _01366_;
  assign _01369_ = sel_oi_one_hot_i[66] & i[34];
  assign _01370_ = sel_oi_one_hot_i[67] & i[50];
  assign _01371_ = _01370_ | _01369_;
  assign _01372_ = _01371_ | _01368_;
  assign _01373_ = sel_oi_one_hot_i[68] & i[66];
  assign _01374_ = sel_oi_one_hot_i[69] & i[82];
  assign _01375_ = _01374_ | _01373_;
  assign _01376_ = sel_oi_one_hot_i[70] & i[98];
  assign _01377_ = sel_oi_one_hot_i[71] & i[114];
  assign _01378_ = _01377_ | _01376_;
  assign _01379_ = _01378_ | _01375_;
  assign _01380_ = _01379_ | _01372_;
  assign _01381_ = sel_oi_one_hot_i[72] & i[130];
  assign _01382_ = sel_oi_one_hot_i[73] & i[146];
  assign _01383_ = _01382_ | _01381_;
  assign _01384_ = sel_oi_one_hot_i[74] & i[162];
  assign _01385_ = sel_oi_one_hot_i[75] & i[178];
  assign _01386_ = _01385_ | _01384_;
  assign _01387_ = _01386_ | _01383_;
  assign _01388_ = sel_oi_one_hot_i[76] & i[194];
  assign _01389_ = sel_oi_one_hot_i[77] & i[210];
  assign _01390_ = _01389_ | _01388_;
  assign _01391_ = sel_oi_one_hot_i[78] & i[226];
  assign _01392_ = sel_oi_one_hot_i[79] & i[242];
  assign _01393_ = _01392_ | _01391_;
  assign _01394_ = _01393_ | _01390_;
  assign _01395_ = _01394_ | _01387_;
  assign o[66] = _01395_ | _01380_;
  assign _01396_ = sel_oi_one_hot_i[64] & i[1];
  assign _01397_ = sel_oi_one_hot_i[65] & i[17];
  assign _01398_ = _01397_ | _01396_;
  assign _01399_ = sel_oi_one_hot_i[66] & i[33];
  assign _01400_ = sel_oi_one_hot_i[67] & i[49];
  assign _01401_ = _01400_ | _01399_;
  assign _01402_ = _01401_ | _01398_;
  assign _01403_ = sel_oi_one_hot_i[68] & i[65];
  assign _01404_ = sel_oi_one_hot_i[69] & i[81];
  assign _01405_ = _01404_ | _01403_;
  assign _01406_ = sel_oi_one_hot_i[70] & i[97];
  assign _01407_ = sel_oi_one_hot_i[71] & i[113];
  assign _01408_ = _01407_ | _01406_;
  assign _01409_ = _01408_ | _01405_;
  assign _01410_ = _01409_ | _01402_;
  assign _01411_ = sel_oi_one_hot_i[72] & i[129];
  assign _01412_ = sel_oi_one_hot_i[73] & i[145];
  assign _01413_ = _01412_ | _01411_;
  assign _01414_ = sel_oi_one_hot_i[74] & i[161];
  assign _01415_ = sel_oi_one_hot_i[75] & i[177];
  assign _01416_ = _01415_ | _01414_;
  assign _01417_ = _01416_ | _01413_;
  assign _01418_ = sel_oi_one_hot_i[76] & i[193];
  assign _01419_ = sel_oi_one_hot_i[77] & i[209];
  assign _01420_ = _01419_ | _01418_;
  assign _01421_ = sel_oi_one_hot_i[78] & i[225];
  assign _01422_ = sel_oi_one_hot_i[79] & i[241];
  assign _01423_ = _01422_ | _01421_;
  assign _01424_ = _01423_ | _01420_;
  assign _01425_ = _01424_ | _01417_;
  assign o[65] = _01425_ | _01410_;
  assign _01426_ = sel_oi_one_hot_i[64] & i[0];
  assign _01427_ = sel_oi_one_hot_i[65] & i[16];
  assign _01428_ = _01427_ | _01426_;
  assign _01429_ = sel_oi_one_hot_i[66] & i[32];
  assign _01430_ = sel_oi_one_hot_i[67] & i[48];
  assign _01431_ = _01430_ | _01429_;
  assign _01432_ = _01431_ | _01428_;
  assign _01433_ = sel_oi_one_hot_i[68] & i[64];
  assign _01434_ = sel_oi_one_hot_i[69] & i[80];
  assign _01435_ = _01434_ | _01433_;
  assign _01436_ = sel_oi_one_hot_i[70] & i[96];
  assign _01437_ = sel_oi_one_hot_i[71] & i[112];
  assign _01438_ = _01437_ | _01436_;
  assign _01439_ = _01438_ | _01435_;
  assign _01440_ = _01439_ | _01432_;
  assign _01441_ = sel_oi_one_hot_i[72] & i[128];
  assign _01442_ = sel_oi_one_hot_i[73] & i[144];
  assign _01443_ = _01442_ | _01441_;
  assign _01444_ = sel_oi_one_hot_i[74] & i[160];
  assign _01445_ = sel_oi_one_hot_i[75] & i[176];
  assign _01446_ = _01445_ | _01444_;
  assign _01447_ = _01446_ | _01443_;
  assign _01448_ = sel_oi_one_hot_i[76] & i[192];
  assign _01449_ = sel_oi_one_hot_i[77] & i[208];
  assign _01450_ = _01449_ | _01448_;
  assign _01451_ = sel_oi_one_hot_i[78] & i[224];
  assign _01452_ = sel_oi_one_hot_i[79] & i[240];
  assign _01453_ = _01452_ | _01451_;
  assign _01454_ = _01453_ | _01450_;
  assign _01455_ = _01454_ | _01447_;
  assign o[64] = _01455_ | _01440_;
  assign _01456_ = sel_oi_one_hot_i[0] & i[7];
  assign _01457_ = sel_oi_one_hot_i[1] & i[23];
  assign _01458_ = _01457_ | _01456_;
  assign _01459_ = sel_oi_one_hot_i[2] & i[39];
  assign _01460_ = sel_oi_one_hot_i[3] & i[55];
  assign _01461_ = _01460_ | _01459_;
  assign _01462_ = _01461_ | _01458_;
  assign _01463_ = sel_oi_one_hot_i[4] & i[71];
  assign _01464_ = sel_oi_one_hot_i[5] & i[87];
  assign _01465_ = _01464_ | _01463_;
  assign _01466_ = sel_oi_one_hot_i[6] & i[103];
  assign _01467_ = sel_oi_one_hot_i[7] & i[119];
  assign _01468_ = _01467_ | _01466_;
  assign _01469_ = _01468_ | _01465_;
  assign _01470_ = _01469_ | _01462_;
  assign _01471_ = sel_oi_one_hot_i[8] & i[135];
  assign _01472_ = sel_oi_one_hot_i[9] & i[151];
  assign _01473_ = _01472_ | _01471_;
  assign _01474_ = sel_oi_one_hot_i[10] & i[167];
  assign _01475_ = sel_oi_one_hot_i[11] & i[183];
  assign _01476_ = _01475_ | _01474_;
  assign _01477_ = _01476_ | _01473_;
  assign _01478_ = sel_oi_one_hot_i[12] & i[199];
  assign _01479_ = sel_oi_one_hot_i[13] & i[215];
  assign _01480_ = _01479_ | _01478_;
  assign _01481_ = sel_oi_one_hot_i[14] & i[231];
  assign _01482_ = sel_oi_one_hot_i[15] & i[247];
  assign _01483_ = _01482_ | _01481_;
  assign _01484_ = _01483_ | _01480_;
  assign _01485_ = _01484_ | _01477_;
  assign o[7] = _01485_ | _01470_;
  assign _01486_ = sel_oi_one_hot_i[80] & i[15];
  assign _01487_ = sel_oi_one_hot_i[81] & i[31];
  assign _01488_ = _01487_ | _01486_;
  assign _01489_ = sel_oi_one_hot_i[82] & i[47];
  assign _01490_ = sel_oi_one_hot_i[83] & i[63];
  assign _01491_ = _01490_ | _01489_;
  assign _01492_ = _01491_ | _01488_;
  assign _01493_ = sel_oi_one_hot_i[84] & i[79];
  assign _01494_ = sel_oi_one_hot_i[85] & i[95];
  assign _01495_ = _01494_ | _01493_;
  assign _01496_ = sel_oi_one_hot_i[86] & i[111];
  assign _01497_ = sel_oi_one_hot_i[87] & i[127];
  assign _01498_ = _01497_ | _01496_;
  assign _01499_ = _01498_ | _01495_;
  assign _01500_ = _01499_ | _01492_;
  assign _01501_ = sel_oi_one_hot_i[88] & i[143];
  assign _01502_ = sel_oi_one_hot_i[89] & i[159];
  assign _01503_ = _01502_ | _01501_;
  assign _01504_ = sel_oi_one_hot_i[90] & i[175];
  assign _01505_ = sel_oi_one_hot_i[91] & i[191];
  assign _01506_ = _01505_ | _01504_;
  assign _01507_ = _01506_ | _01503_;
  assign _01508_ = sel_oi_one_hot_i[92] & i[207];
  assign _01509_ = sel_oi_one_hot_i[93] & i[223];
  assign _01510_ = _01509_ | _01508_;
  assign _01511_ = sel_oi_one_hot_i[94] & i[239];
  assign _01512_ = sel_oi_one_hot_i[95] & i[255];
  assign _01513_ = _01512_ | _01511_;
  assign _01514_ = _01513_ | _01510_;
  assign _01515_ = _01514_ | _01507_;
  assign o[95] = _01515_ | _01500_;
  assign _01516_ = sel_oi_one_hot_i[80] & i[14];
  assign _01517_ = sel_oi_one_hot_i[81] & i[30];
  assign _01518_ = _01517_ | _01516_;
  assign _01519_ = sel_oi_one_hot_i[82] & i[46];
  assign _01520_ = sel_oi_one_hot_i[83] & i[62];
  assign _01521_ = _01520_ | _01519_;
  assign _01522_ = _01521_ | _01518_;
  assign _01523_ = sel_oi_one_hot_i[84] & i[78];
  assign _01524_ = sel_oi_one_hot_i[85] & i[94];
  assign _01525_ = _01524_ | _01523_;
  assign _01526_ = sel_oi_one_hot_i[86] & i[110];
  assign _01527_ = sel_oi_one_hot_i[87] & i[126];
  assign _01528_ = _01527_ | _01526_;
  assign _01529_ = _01528_ | _01525_;
  assign _01530_ = _01529_ | _01522_;
  assign _01531_ = sel_oi_one_hot_i[88] & i[142];
  assign _01532_ = sel_oi_one_hot_i[89] & i[158];
  assign _01533_ = _01532_ | _01531_;
  assign _01534_ = sel_oi_one_hot_i[90] & i[174];
  assign _01535_ = sel_oi_one_hot_i[91] & i[190];
  assign _01536_ = _01535_ | _01534_;
  assign _01537_ = _01536_ | _01533_;
  assign _01538_ = sel_oi_one_hot_i[92] & i[206];
  assign _01539_ = sel_oi_one_hot_i[93] & i[222];
  assign _01540_ = _01539_ | _01538_;
  assign _01541_ = sel_oi_one_hot_i[94] & i[238];
  assign _01542_ = sel_oi_one_hot_i[95] & i[254];
  assign _01543_ = _01542_ | _01541_;
  assign _01544_ = _01543_ | _01540_;
  assign _01545_ = _01544_ | _01537_;
  assign o[94] = _01545_ | _01530_;
  assign _01546_ = sel_oi_one_hot_i[80] & i[13];
  assign _01547_ = sel_oi_one_hot_i[81] & i[29];
  assign _01548_ = _01547_ | _01546_;
  assign _01549_ = sel_oi_one_hot_i[82] & i[45];
  assign _01550_ = sel_oi_one_hot_i[83] & i[61];
  assign _01551_ = _01550_ | _01549_;
  assign _01552_ = _01551_ | _01548_;
  assign _01553_ = sel_oi_one_hot_i[84] & i[77];
  assign _01554_ = sel_oi_one_hot_i[85] & i[93];
  assign _01555_ = _01554_ | _01553_;
  assign _01556_ = sel_oi_one_hot_i[86] & i[109];
  assign _01557_ = sel_oi_one_hot_i[87] & i[125];
  assign _01558_ = _01557_ | _01556_;
  assign _01559_ = _01558_ | _01555_;
  assign _01560_ = _01559_ | _01552_;
  assign _01561_ = sel_oi_one_hot_i[88] & i[141];
  assign _01562_ = sel_oi_one_hot_i[89] & i[157];
  assign _01563_ = _01562_ | _01561_;
  assign _01564_ = sel_oi_one_hot_i[90] & i[173];
  assign _01565_ = sel_oi_one_hot_i[91] & i[189];
  assign _01566_ = _01565_ | _01564_;
  assign _01567_ = _01566_ | _01563_;
  assign _01568_ = sel_oi_one_hot_i[92] & i[205];
  assign _01569_ = sel_oi_one_hot_i[93] & i[221];
  assign _01570_ = _01569_ | _01568_;
  assign _01571_ = sel_oi_one_hot_i[94] & i[237];
  assign _01572_ = sel_oi_one_hot_i[95] & i[253];
  assign _01573_ = _01572_ | _01571_;
  assign _01574_ = _01573_ | _01570_;
  assign _01575_ = _01574_ | _01567_;
  assign o[93] = _01575_ | _01560_;
  assign _01576_ = sel_oi_one_hot_i[80] & i[12];
  assign _01577_ = sel_oi_one_hot_i[81] & i[28];
  assign _01578_ = _01577_ | _01576_;
  assign _01579_ = sel_oi_one_hot_i[82] & i[44];
  assign _01580_ = sel_oi_one_hot_i[83] & i[60];
  assign _01581_ = _01580_ | _01579_;
  assign _01582_ = _01581_ | _01578_;
  assign _01583_ = sel_oi_one_hot_i[84] & i[76];
  assign _01584_ = sel_oi_one_hot_i[85] & i[92];
  assign _01585_ = _01584_ | _01583_;
  assign _01586_ = sel_oi_one_hot_i[86] & i[108];
  assign _01587_ = sel_oi_one_hot_i[87] & i[124];
  assign _01588_ = _01587_ | _01586_;
  assign _01589_ = _01588_ | _01585_;
  assign _01590_ = _01589_ | _01582_;
  assign _01591_ = sel_oi_one_hot_i[88] & i[140];
  assign _01592_ = sel_oi_one_hot_i[89] & i[156];
  assign _01593_ = _01592_ | _01591_;
  assign _01594_ = sel_oi_one_hot_i[90] & i[172];
  assign _01595_ = sel_oi_one_hot_i[91] & i[188];
  assign _01596_ = _01595_ | _01594_;
  assign _01597_ = _01596_ | _01593_;
  assign _01598_ = sel_oi_one_hot_i[92] & i[204];
  assign _01599_ = sel_oi_one_hot_i[93] & i[220];
  assign _01600_ = _01599_ | _01598_;
  assign _01601_ = sel_oi_one_hot_i[94] & i[236];
  assign _01602_ = sel_oi_one_hot_i[95] & i[252];
  assign _01603_ = _01602_ | _01601_;
  assign _01604_ = _01603_ | _01600_;
  assign _01605_ = _01604_ | _01597_;
  assign o[92] = _01605_ | _01590_;
  assign _01606_ = sel_oi_one_hot_i[0] & i[6];
  assign _01607_ = sel_oi_one_hot_i[1] & i[22];
  assign _01608_ = _01607_ | _01606_;
  assign _01609_ = sel_oi_one_hot_i[2] & i[38];
  assign _01610_ = sel_oi_one_hot_i[3] & i[54];
  assign _01611_ = _01610_ | _01609_;
  assign _01612_ = _01611_ | _01608_;
  assign _01613_ = sel_oi_one_hot_i[4] & i[70];
  assign _01614_ = sel_oi_one_hot_i[5] & i[86];
  assign _01615_ = _01614_ | _01613_;
  assign _01616_ = sel_oi_one_hot_i[6] & i[102];
  assign _01617_ = sel_oi_one_hot_i[7] & i[118];
  assign _01618_ = _01617_ | _01616_;
  assign _01619_ = _01618_ | _01615_;
  assign _01620_ = _01619_ | _01612_;
  assign _01621_ = sel_oi_one_hot_i[8] & i[134];
  assign _01622_ = sel_oi_one_hot_i[9] & i[150];
  assign _01623_ = _01622_ | _01621_;
  assign _01624_ = sel_oi_one_hot_i[10] & i[166];
  assign _01625_ = sel_oi_one_hot_i[11] & i[182];
  assign _01626_ = _01625_ | _01624_;
  assign _01627_ = _01626_ | _01623_;
  assign _01628_ = sel_oi_one_hot_i[12] & i[198];
  assign _01629_ = sel_oi_one_hot_i[13] & i[214];
  assign _01630_ = _01629_ | _01628_;
  assign _01631_ = sel_oi_one_hot_i[14] & i[230];
  assign _01632_ = sel_oi_one_hot_i[15] & i[246];
  assign _01633_ = _01632_ | _01631_;
  assign _01634_ = _01633_ | _01630_;
  assign _01635_ = _01634_ | _01627_;
  assign o[6] = _01635_ | _01620_;
  assign _01636_ = sel_oi_one_hot_i[80] & i[11];
  assign _01637_ = sel_oi_one_hot_i[81] & i[27];
  assign _01638_ = _01637_ | _01636_;
  assign _01639_ = sel_oi_one_hot_i[82] & i[43];
  assign _01640_ = sel_oi_one_hot_i[83] & i[59];
  assign _01641_ = _01640_ | _01639_;
  assign _01642_ = _01641_ | _01638_;
  assign _01643_ = sel_oi_one_hot_i[84] & i[75];
  assign _01644_ = sel_oi_one_hot_i[85] & i[91];
  assign _01645_ = _01644_ | _01643_;
  assign _01646_ = sel_oi_one_hot_i[86] & i[107];
  assign _01647_ = sel_oi_one_hot_i[87] & i[123];
  assign _01648_ = _01647_ | _01646_;
  assign _01649_ = _01648_ | _01645_;
  assign _01650_ = _01649_ | _01642_;
  assign _01651_ = sel_oi_one_hot_i[88] & i[139];
  assign _01652_ = sel_oi_one_hot_i[89] & i[155];
  assign _01653_ = _01652_ | _01651_;
  assign _01654_ = sel_oi_one_hot_i[90] & i[171];
  assign _01655_ = sel_oi_one_hot_i[91] & i[187];
  assign _01656_ = _01655_ | _01654_;
  assign _01657_ = _01656_ | _01653_;
  assign _01658_ = sel_oi_one_hot_i[92] & i[203];
  assign _01659_ = sel_oi_one_hot_i[93] & i[219];
  assign _01660_ = _01659_ | _01658_;
  assign _01661_ = sel_oi_one_hot_i[94] & i[235];
  assign _01662_ = sel_oi_one_hot_i[95] & i[251];
  assign _01663_ = _01662_ | _01661_;
  assign _01664_ = _01663_ | _01660_;
  assign _01665_ = _01664_ | _01657_;
  assign o[91] = _01665_ | _01650_;
  assign _01666_ = sel_oi_one_hot_i[80] & i[10];
  assign _01667_ = sel_oi_one_hot_i[81] & i[26];
  assign _01668_ = _01667_ | _01666_;
  assign _01669_ = sel_oi_one_hot_i[82] & i[42];
  assign _01670_ = sel_oi_one_hot_i[83] & i[58];
  assign _01671_ = _01670_ | _01669_;
  assign _01672_ = _01671_ | _01668_;
  assign _01673_ = sel_oi_one_hot_i[84] & i[74];
  assign _01674_ = sel_oi_one_hot_i[85] & i[90];
  assign _01675_ = _01674_ | _01673_;
  assign _01676_ = sel_oi_one_hot_i[86] & i[106];
  assign _01677_ = sel_oi_one_hot_i[87] & i[122];
  assign _01678_ = _01677_ | _01676_;
  assign _01679_ = _01678_ | _01675_;
  assign _01680_ = _01679_ | _01672_;
  assign _01681_ = sel_oi_one_hot_i[88] & i[138];
  assign _01682_ = sel_oi_one_hot_i[89] & i[154];
  assign _01683_ = _01682_ | _01681_;
  assign _01684_ = sel_oi_one_hot_i[90] & i[170];
  assign _01685_ = sel_oi_one_hot_i[91] & i[186];
  assign _01686_ = _01685_ | _01684_;
  assign _01687_ = _01686_ | _01683_;
  assign _01688_ = sel_oi_one_hot_i[92] & i[202];
  assign _01689_ = sel_oi_one_hot_i[93] & i[218];
  assign _01690_ = _01689_ | _01688_;
  assign _01691_ = sel_oi_one_hot_i[94] & i[234];
  assign _01692_ = sel_oi_one_hot_i[95] & i[250];
  assign _01693_ = _01692_ | _01691_;
  assign _01694_ = _01693_ | _01690_;
  assign _01695_ = _01694_ | _01687_;
  assign o[90] = _01695_ | _01680_;
  assign _01696_ = sel_oi_one_hot_i[80] & i[9];
  assign _01697_ = sel_oi_one_hot_i[81] & i[25];
  assign _01698_ = _01697_ | _01696_;
  assign _01699_ = sel_oi_one_hot_i[82] & i[41];
  assign _01700_ = sel_oi_one_hot_i[83] & i[57];
  assign _01701_ = _01700_ | _01699_;
  assign _01702_ = _01701_ | _01698_;
  assign _01703_ = sel_oi_one_hot_i[84] & i[73];
  assign _01704_ = sel_oi_one_hot_i[85] & i[89];
  assign _01705_ = _01704_ | _01703_;
  assign _01706_ = sel_oi_one_hot_i[86] & i[105];
  assign _01707_ = sel_oi_one_hot_i[87] & i[121];
  assign _01708_ = _01707_ | _01706_;
  assign _01709_ = _01708_ | _01705_;
  assign _01710_ = _01709_ | _01702_;
  assign _01711_ = sel_oi_one_hot_i[88] & i[137];
  assign _01712_ = sel_oi_one_hot_i[89] & i[153];
  assign _01713_ = _01712_ | _01711_;
  assign _01714_ = sel_oi_one_hot_i[90] & i[169];
  assign _01715_ = sel_oi_one_hot_i[91] & i[185];
  assign _01716_ = _01715_ | _01714_;
  assign _01717_ = _01716_ | _01713_;
  assign _01718_ = sel_oi_one_hot_i[92] & i[201];
  assign _01719_ = sel_oi_one_hot_i[93] & i[217];
  assign _01720_ = _01719_ | _01718_;
  assign _01721_ = sel_oi_one_hot_i[94] & i[233];
  assign _01722_ = sel_oi_one_hot_i[95] & i[249];
  assign _01723_ = _01722_ | _01721_;
  assign _01724_ = _01723_ | _01720_;
  assign _01725_ = _01724_ | _01717_;
  assign o[89] = _01725_ | _01710_;
  assign _01726_ = sel_oi_one_hot_i[80] & i[8];
  assign _01727_ = sel_oi_one_hot_i[81] & i[24];
  assign _01728_ = _01727_ | _01726_;
  assign _01729_ = sel_oi_one_hot_i[82] & i[40];
  assign _01730_ = sel_oi_one_hot_i[83] & i[56];
  assign _01731_ = _01730_ | _01729_;
  assign _01732_ = _01731_ | _01728_;
  assign _01733_ = sel_oi_one_hot_i[84] & i[72];
  assign _01734_ = sel_oi_one_hot_i[85] & i[88];
  assign _01735_ = _01734_ | _01733_;
  assign _01736_ = sel_oi_one_hot_i[86] & i[104];
  assign _01737_ = sel_oi_one_hot_i[87] & i[120];
  assign _01738_ = _01737_ | _01736_;
  assign _01739_ = _01738_ | _01735_;
  assign _01740_ = _01739_ | _01732_;
  assign _01741_ = sel_oi_one_hot_i[88] & i[136];
  assign _01742_ = sel_oi_one_hot_i[89] & i[152];
  assign _01743_ = _01742_ | _01741_;
  assign _01744_ = sel_oi_one_hot_i[90] & i[168];
  assign _01745_ = sel_oi_one_hot_i[91] & i[184];
  assign _01746_ = _01745_ | _01744_;
  assign _01747_ = _01746_ | _01743_;
  assign _01748_ = sel_oi_one_hot_i[92] & i[200];
  assign _01749_ = sel_oi_one_hot_i[93] & i[216];
  assign _01750_ = _01749_ | _01748_;
  assign _01751_ = sel_oi_one_hot_i[94] & i[232];
  assign _01752_ = sel_oi_one_hot_i[95] & i[248];
  assign _01753_ = _01752_ | _01751_;
  assign _01754_ = _01753_ | _01750_;
  assign _01755_ = _01754_ | _01747_;
  assign o[88] = _01755_ | _01740_;
  assign _01756_ = sel_oi_one_hot_i[80] & i[7];
  assign _01757_ = sel_oi_one_hot_i[81] & i[23];
  assign _01758_ = _01757_ | _01756_;
  assign _01759_ = sel_oi_one_hot_i[82] & i[39];
  assign _01760_ = sel_oi_one_hot_i[83] & i[55];
  assign _01761_ = _01760_ | _01759_;
  assign _01762_ = _01761_ | _01758_;
  assign _01763_ = sel_oi_one_hot_i[84] & i[71];
  assign _01764_ = sel_oi_one_hot_i[85] & i[87];
  assign _01765_ = _01764_ | _01763_;
  assign _01766_ = sel_oi_one_hot_i[86] & i[103];
  assign _01767_ = sel_oi_one_hot_i[87] & i[119];
  assign _01768_ = _01767_ | _01766_;
  assign _01769_ = _01768_ | _01765_;
  assign _01770_ = _01769_ | _01762_;
  assign _01771_ = sel_oi_one_hot_i[88] & i[135];
  assign _01772_ = sel_oi_one_hot_i[89] & i[151];
  assign _01773_ = _01772_ | _01771_;
  assign _01774_ = sel_oi_one_hot_i[90] & i[167];
  assign _01775_ = sel_oi_one_hot_i[91] & i[183];
  assign _01776_ = _01775_ | _01774_;
  assign _01777_ = _01776_ | _01773_;
  assign _01778_ = sel_oi_one_hot_i[92] & i[199];
  assign _01779_ = sel_oi_one_hot_i[93] & i[215];
  assign _01780_ = _01779_ | _01778_;
  assign _01781_ = sel_oi_one_hot_i[94] & i[231];
  assign _01782_ = sel_oi_one_hot_i[95] & i[247];
  assign _01783_ = _01782_ | _01781_;
  assign _01784_ = _01783_ | _01780_;
  assign _01785_ = _01784_ | _01777_;
  assign o[87] = _01785_ | _01770_;
  assign _01786_ = sel_oi_one_hot_i[80] & i[6];
  assign _01787_ = sel_oi_one_hot_i[81] & i[22];
  assign _01788_ = _01787_ | _01786_;
  assign _01789_ = sel_oi_one_hot_i[82] & i[38];
  assign _01790_ = sel_oi_one_hot_i[83] & i[54];
  assign _01791_ = _01790_ | _01789_;
  assign _01792_ = _01791_ | _01788_;
  assign _01793_ = sel_oi_one_hot_i[84] & i[70];
  assign _01794_ = sel_oi_one_hot_i[85] & i[86];
  assign _01795_ = _01794_ | _01793_;
  assign _01796_ = sel_oi_one_hot_i[86] & i[102];
  assign _01797_ = sel_oi_one_hot_i[87] & i[118];
  assign _01798_ = _01797_ | _01796_;
  assign _01799_ = _01798_ | _01795_;
  assign _01800_ = _01799_ | _01792_;
  assign _01801_ = sel_oi_one_hot_i[88] & i[134];
  assign _01802_ = sel_oi_one_hot_i[89] & i[150];
  assign _01803_ = _01802_ | _01801_;
  assign _01804_ = sel_oi_one_hot_i[90] & i[166];
  assign _01805_ = sel_oi_one_hot_i[91] & i[182];
  assign _01806_ = _01805_ | _01804_;
  assign _01807_ = _01806_ | _01803_;
  assign _01808_ = sel_oi_one_hot_i[92] & i[198];
  assign _01809_ = sel_oi_one_hot_i[93] & i[214];
  assign _01810_ = _01809_ | _01808_;
  assign _01811_ = sel_oi_one_hot_i[94] & i[230];
  assign _01812_ = sel_oi_one_hot_i[95] & i[246];
  assign _01813_ = _01812_ | _01811_;
  assign _01814_ = _01813_ | _01810_;
  assign _01815_ = _01814_ | _01807_;
  assign o[86] = _01815_ | _01800_;
  assign _01816_ = sel_oi_one_hot_i[80] & i[5];
  assign _01817_ = sel_oi_one_hot_i[81] & i[21];
  assign _01818_ = _01817_ | _01816_;
  assign _01819_ = sel_oi_one_hot_i[82] & i[37];
  assign _01820_ = sel_oi_one_hot_i[83] & i[53];
  assign _01821_ = _01820_ | _01819_;
  assign _01822_ = _01821_ | _01818_;
  assign _01823_ = sel_oi_one_hot_i[84] & i[69];
  assign _01824_ = sel_oi_one_hot_i[85] & i[85];
  assign _01825_ = _01824_ | _01823_;
  assign _01826_ = sel_oi_one_hot_i[86] & i[101];
  assign _01827_ = sel_oi_one_hot_i[87] & i[117];
  assign _01828_ = _01827_ | _01826_;
  assign _01829_ = _01828_ | _01825_;
  assign _01830_ = _01829_ | _01822_;
  assign _01831_ = sel_oi_one_hot_i[88] & i[133];
  assign _01832_ = sel_oi_one_hot_i[89] & i[149];
  assign _01833_ = _01832_ | _01831_;
  assign _01834_ = sel_oi_one_hot_i[90] & i[165];
  assign _01835_ = sel_oi_one_hot_i[91] & i[181];
  assign _01836_ = _01835_ | _01834_;
  assign _01837_ = _01836_ | _01833_;
  assign _01838_ = sel_oi_one_hot_i[92] & i[197];
  assign _01839_ = sel_oi_one_hot_i[93] & i[213];
  assign _01840_ = _01839_ | _01838_;
  assign _01841_ = sel_oi_one_hot_i[94] & i[229];
  assign _01842_ = sel_oi_one_hot_i[95] & i[245];
  assign _01843_ = _01842_ | _01841_;
  assign _01844_ = _01843_ | _01840_;
  assign _01845_ = _01844_ | _01837_;
  assign o[85] = _01845_ | _01830_;
  assign _01846_ = sel_oi_one_hot_i[80] & i[4];
  assign _01847_ = sel_oi_one_hot_i[81] & i[20];
  assign _01848_ = _01847_ | _01846_;
  assign _01849_ = sel_oi_one_hot_i[82] & i[36];
  assign _01850_ = sel_oi_one_hot_i[83] & i[52];
  assign _01851_ = _01850_ | _01849_;
  assign _01852_ = _01851_ | _01848_;
  assign _01853_ = sel_oi_one_hot_i[84] & i[68];
  assign _01854_ = sel_oi_one_hot_i[85] & i[84];
  assign _01855_ = _01854_ | _01853_;
  assign _01856_ = sel_oi_one_hot_i[86] & i[100];
  assign _01857_ = sel_oi_one_hot_i[87] & i[116];
  assign _01858_ = _01857_ | _01856_;
  assign _01859_ = _01858_ | _01855_;
  assign _01860_ = _01859_ | _01852_;
  assign _01861_ = sel_oi_one_hot_i[88] & i[132];
  assign _01862_ = sel_oi_one_hot_i[89] & i[148];
  assign _01863_ = _01862_ | _01861_;
  assign _01864_ = sel_oi_one_hot_i[90] & i[164];
  assign _01865_ = sel_oi_one_hot_i[91] & i[180];
  assign _01866_ = _01865_ | _01864_;
  assign _01867_ = _01866_ | _01863_;
  assign _01868_ = sel_oi_one_hot_i[92] & i[196];
  assign _01869_ = sel_oi_one_hot_i[93] & i[212];
  assign _01870_ = _01869_ | _01868_;
  assign _01871_ = sel_oi_one_hot_i[94] & i[228];
  assign _01872_ = sel_oi_one_hot_i[95] & i[244];
  assign _01873_ = _01872_ | _01871_;
  assign _01874_ = _01873_ | _01870_;
  assign _01875_ = _01874_ | _01867_;
  assign o[84] = _01875_ | _01860_;
  assign _01876_ = sel_oi_one_hot_i[80] & i[3];
  assign _01877_ = sel_oi_one_hot_i[81] & i[19];
  assign _01878_ = _01877_ | _01876_;
  assign _01879_ = sel_oi_one_hot_i[82] & i[35];
  assign _01880_ = sel_oi_one_hot_i[83] & i[51];
  assign _01881_ = _01880_ | _01879_;
  assign _01882_ = _01881_ | _01878_;
  assign _01883_ = sel_oi_one_hot_i[84] & i[67];
  assign _01884_ = sel_oi_one_hot_i[85] & i[83];
  assign _01885_ = _01884_ | _01883_;
  assign _01886_ = sel_oi_one_hot_i[86] & i[99];
  assign _01887_ = sel_oi_one_hot_i[87] & i[115];
  assign _01888_ = _01887_ | _01886_;
  assign _01889_ = _01888_ | _01885_;
  assign _01890_ = _01889_ | _01882_;
  assign _01891_ = sel_oi_one_hot_i[88] & i[131];
  assign _01892_ = sel_oi_one_hot_i[89] & i[147];
  assign _01893_ = _01892_ | _01891_;
  assign _01894_ = sel_oi_one_hot_i[90] & i[163];
  assign _01895_ = sel_oi_one_hot_i[91] & i[179];
  assign _01896_ = _01895_ | _01894_;
  assign _01897_ = _01896_ | _01893_;
  assign _01898_ = sel_oi_one_hot_i[92] & i[195];
  assign _01899_ = sel_oi_one_hot_i[93] & i[211];
  assign _01900_ = _01899_ | _01898_;
  assign _01901_ = sel_oi_one_hot_i[94] & i[227];
  assign _01902_ = sel_oi_one_hot_i[95] & i[243];
  assign _01903_ = _01902_ | _01901_;
  assign _01904_ = _01903_ | _01900_;
  assign _01905_ = _01904_ | _01897_;
  assign o[83] = _01905_ | _01890_;
  assign _01906_ = sel_oi_one_hot_i[80] & i[2];
  assign _01907_ = sel_oi_one_hot_i[81] & i[18];
  assign _01908_ = _01907_ | _01906_;
  assign _01909_ = sel_oi_one_hot_i[82] & i[34];
  assign _01910_ = sel_oi_one_hot_i[83] & i[50];
  assign _01911_ = _01910_ | _01909_;
  assign _01912_ = _01911_ | _01908_;
  assign _01913_ = sel_oi_one_hot_i[84] & i[66];
  assign _01914_ = sel_oi_one_hot_i[85] & i[82];
  assign _01915_ = _01914_ | _01913_;
  assign _01916_ = sel_oi_one_hot_i[86] & i[98];
  assign _01917_ = sel_oi_one_hot_i[87] & i[114];
  assign _01918_ = _01917_ | _01916_;
  assign _01919_ = _01918_ | _01915_;
  assign _01920_ = _01919_ | _01912_;
  assign _01921_ = sel_oi_one_hot_i[88] & i[130];
  assign _01922_ = sel_oi_one_hot_i[89] & i[146];
  assign _01923_ = _01922_ | _01921_;
  assign _01924_ = sel_oi_one_hot_i[90] & i[162];
  assign _01925_ = sel_oi_one_hot_i[91] & i[178];
  assign _01926_ = _01925_ | _01924_;
  assign _01927_ = _01926_ | _01923_;
  assign _01928_ = sel_oi_one_hot_i[92] & i[194];
  assign _01929_ = sel_oi_one_hot_i[93] & i[210];
  assign _01930_ = _01929_ | _01928_;
  assign _01931_ = sel_oi_one_hot_i[94] & i[226];
  assign _01932_ = sel_oi_one_hot_i[95] & i[242];
  assign _01933_ = _01932_ | _01931_;
  assign _01934_ = _01933_ | _01930_;
  assign _01935_ = _01934_ | _01927_;
  assign o[82] = _01935_ | _01920_;
  assign _01936_ = sel_oi_one_hot_i[0] & i[5];
  assign _01937_ = sel_oi_one_hot_i[1] & i[21];
  assign _01938_ = _01937_ | _01936_;
  assign _01939_ = sel_oi_one_hot_i[2] & i[37];
  assign _01940_ = sel_oi_one_hot_i[3] & i[53];
  assign _01941_ = _01940_ | _01939_;
  assign _01942_ = _01941_ | _01938_;
  assign _01943_ = sel_oi_one_hot_i[4] & i[69];
  assign _01944_ = sel_oi_one_hot_i[5] & i[85];
  assign _01945_ = _01944_ | _01943_;
  assign _01946_ = sel_oi_one_hot_i[6] & i[101];
  assign _01947_ = sel_oi_one_hot_i[7] & i[117];
  assign _01948_ = _01947_ | _01946_;
  assign _01949_ = _01948_ | _01945_;
  assign _01950_ = _01949_ | _01942_;
  assign _01951_ = sel_oi_one_hot_i[8] & i[133];
  assign _01952_ = sel_oi_one_hot_i[9] & i[149];
  assign _01953_ = _01952_ | _01951_;
  assign _01954_ = sel_oi_one_hot_i[10] & i[165];
  assign _01955_ = sel_oi_one_hot_i[11] & i[181];
  assign _01956_ = _01955_ | _01954_;
  assign _01957_ = _01956_ | _01953_;
  assign _01958_ = sel_oi_one_hot_i[12] & i[197];
  assign _01959_ = sel_oi_one_hot_i[13] & i[213];
  assign _01960_ = _01959_ | _01958_;
  assign _01961_ = sel_oi_one_hot_i[14] & i[229];
  assign _01962_ = sel_oi_one_hot_i[15] & i[245];
  assign _01963_ = _01962_ | _01961_;
  assign _01964_ = _01963_ | _01960_;
  assign _01965_ = _01964_ | _01957_;
  assign o[5] = _01965_ | _01950_;
  assign _01966_ = sel_oi_one_hot_i[80] & i[1];
  assign _01967_ = sel_oi_one_hot_i[81] & i[17];
  assign _01968_ = _01967_ | _01966_;
  assign _01969_ = sel_oi_one_hot_i[82] & i[33];
  assign _01970_ = sel_oi_one_hot_i[83] & i[49];
  assign _01971_ = _01970_ | _01969_;
  assign _01972_ = _01971_ | _01968_;
  assign _01973_ = sel_oi_one_hot_i[84] & i[65];
  assign _01974_ = sel_oi_one_hot_i[85] & i[81];
  assign _01975_ = _01974_ | _01973_;
  assign _01976_ = sel_oi_one_hot_i[86] & i[97];
  assign _01977_ = sel_oi_one_hot_i[87] & i[113];
  assign _01978_ = _01977_ | _01976_;
  assign _01979_ = _01978_ | _01975_;
  assign _01980_ = _01979_ | _01972_;
  assign _01981_ = sel_oi_one_hot_i[88] & i[129];
  assign _01982_ = sel_oi_one_hot_i[89] & i[145];
  assign _01983_ = _01982_ | _01981_;
  assign _01984_ = sel_oi_one_hot_i[90] & i[161];
  assign _01985_ = sel_oi_one_hot_i[91] & i[177];
  assign _01986_ = _01985_ | _01984_;
  assign _01987_ = _01986_ | _01983_;
  assign _01988_ = sel_oi_one_hot_i[92] & i[193];
  assign _01989_ = sel_oi_one_hot_i[93] & i[209];
  assign _01990_ = _01989_ | _01988_;
  assign _01991_ = sel_oi_one_hot_i[94] & i[225];
  assign _01992_ = sel_oi_one_hot_i[95] & i[241];
  assign _01993_ = _01992_ | _01991_;
  assign _01994_ = _01993_ | _01990_;
  assign _01995_ = _01994_ | _01987_;
  assign o[81] = _01995_ | _01980_;
  assign _01996_ = sel_oi_one_hot_i[80] & i[0];
  assign _01997_ = sel_oi_one_hot_i[81] & i[16];
  assign _01998_ = _01997_ | _01996_;
  assign _01999_ = sel_oi_one_hot_i[82] & i[32];
  assign _02000_ = sel_oi_one_hot_i[83] & i[48];
  assign _02001_ = _02000_ | _01999_;
  assign _02002_ = _02001_ | _01998_;
  assign _02003_ = sel_oi_one_hot_i[84] & i[64];
  assign _02004_ = sel_oi_one_hot_i[85] & i[80];
  assign _02005_ = _02004_ | _02003_;
  assign _02006_ = sel_oi_one_hot_i[86] & i[96];
  assign _02007_ = sel_oi_one_hot_i[87] & i[112];
  assign _02008_ = _02007_ | _02006_;
  assign _02009_ = _02008_ | _02005_;
  assign _02010_ = _02009_ | _02002_;
  assign _02011_ = sel_oi_one_hot_i[88] & i[128];
  assign _02012_ = sel_oi_one_hot_i[89] & i[144];
  assign _02013_ = _02012_ | _02011_;
  assign _02014_ = sel_oi_one_hot_i[90] & i[160];
  assign _02015_ = sel_oi_one_hot_i[91] & i[176];
  assign _02016_ = _02015_ | _02014_;
  assign _02017_ = _02016_ | _02013_;
  assign _02018_ = sel_oi_one_hot_i[92] & i[192];
  assign _02019_ = sel_oi_one_hot_i[93] & i[208];
  assign _02020_ = _02019_ | _02018_;
  assign _02021_ = sel_oi_one_hot_i[94] & i[224];
  assign _02022_ = sel_oi_one_hot_i[95] & i[240];
  assign _02023_ = _02022_ | _02021_;
  assign _02024_ = _02023_ | _02020_;
  assign _02025_ = _02024_ | _02017_;
  assign o[80] = _02025_ | _02010_;
  assign _02026_ = sel_oi_one_hot_i[0] & i[4];
  assign _02027_ = sel_oi_one_hot_i[1] & i[20];
  assign _02028_ = _02027_ | _02026_;
  assign _02029_ = sel_oi_one_hot_i[2] & i[36];
  assign _02030_ = sel_oi_one_hot_i[3] & i[52];
  assign _02031_ = _02030_ | _02029_;
  assign _02032_ = _02031_ | _02028_;
  assign _02033_ = sel_oi_one_hot_i[4] & i[68];
  assign _02034_ = sel_oi_one_hot_i[5] & i[84];
  assign _02035_ = _02034_ | _02033_;
  assign _02036_ = sel_oi_one_hot_i[6] & i[100];
  assign _02037_ = sel_oi_one_hot_i[7] & i[116];
  assign _02038_ = _02037_ | _02036_;
  assign _02039_ = _02038_ | _02035_;
  assign _02040_ = _02039_ | _02032_;
  assign _02041_ = sel_oi_one_hot_i[8] & i[132];
  assign _02042_ = sel_oi_one_hot_i[9] & i[148];
  assign _02043_ = _02042_ | _02041_;
  assign _02044_ = sel_oi_one_hot_i[10] & i[164];
  assign _02045_ = sel_oi_one_hot_i[11] & i[180];
  assign _02046_ = _02045_ | _02044_;
  assign _02047_ = _02046_ | _02043_;
  assign _02048_ = sel_oi_one_hot_i[12] & i[196];
  assign _02049_ = sel_oi_one_hot_i[13] & i[212];
  assign _02050_ = _02049_ | _02048_;
  assign _02051_ = sel_oi_one_hot_i[14] & i[228];
  assign _02052_ = sel_oi_one_hot_i[15] & i[244];
  assign _02053_ = _02052_ | _02051_;
  assign _02054_ = _02053_ | _02050_;
  assign _02055_ = _02054_ | _02047_;
  assign o[4] = _02055_ | _02040_;
  assign _02056_ = sel_oi_one_hot_i[96] & i[15];
  assign _02057_ = sel_oi_one_hot_i[97] & i[31];
  assign _02058_ = _02057_ | _02056_;
  assign _02059_ = sel_oi_one_hot_i[98] & i[47];
  assign _02060_ = sel_oi_one_hot_i[99] & i[63];
  assign _02061_ = _02060_ | _02059_;
  assign _02062_ = _02061_ | _02058_;
  assign _02063_ = sel_oi_one_hot_i[100] & i[79];
  assign _02064_ = sel_oi_one_hot_i[101] & i[95];
  assign _02065_ = _02064_ | _02063_;
  assign _02066_ = sel_oi_one_hot_i[102] & i[111];
  assign _02067_ = sel_oi_one_hot_i[103] & i[127];
  assign _02068_ = _02067_ | _02066_;
  assign _02069_ = _02068_ | _02065_;
  assign _02070_ = _02069_ | _02062_;
  assign _02071_ = sel_oi_one_hot_i[104] & i[143];
  assign _02072_ = sel_oi_one_hot_i[105] & i[159];
  assign _02073_ = _02072_ | _02071_;
  assign _02074_ = sel_oi_one_hot_i[106] & i[175];
  assign _02075_ = sel_oi_one_hot_i[107] & i[191];
  assign _02076_ = _02075_ | _02074_;
  assign _02077_ = _02076_ | _02073_;
  assign _02078_ = sel_oi_one_hot_i[108] & i[207];
  assign _02079_ = sel_oi_one_hot_i[109] & i[223];
  assign _02080_ = _02079_ | _02078_;
  assign _02081_ = sel_oi_one_hot_i[110] & i[239];
  assign _02082_ = sel_oi_one_hot_i[111] & i[255];
  assign _02083_ = _02082_ | _02081_;
  assign _02084_ = _02083_ | _02080_;
  assign _02085_ = _02084_ | _02077_;
  assign o[111] = _02085_ | _02070_;
  assign _02086_ = sel_oi_one_hot_i[96] & i[14];
  assign _02087_ = sel_oi_one_hot_i[97] & i[30];
  assign _02088_ = _02087_ | _02086_;
  assign _02089_ = sel_oi_one_hot_i[98] & i[46];
  assign _02090_ = sel_oi_one_hot_i[99] & i[62];
  assign _02091_ = _02090_ | _02089_;
  assign _02092_ = _02091_ | _02088_;
  assign _02093_ = sel_oi_one_hot_i[100] & i[78];
  assign _02094_ = sel_oi_one_hot_i[101] & i[94];
  assign _02095_ = _02094_ | _02093_;
  assign _02096_ = sel_oi_one_hot_i[102] & i[110];
  assign _02097_ = sel_oi_one_hot_i[103] & i[126];
  assign _02098_ = _02097_ | _02096_;
  assign _02099_ = _02098_ | _02095_;
  assign _02100_ = _02099_ | _02092_;
  assign _02101_ = sel_oi_one_hot_i[104] & i[142];
  assign _02102_ = sel_oi_one_hot_i[105] & i[158];
  assign _02103_ = _02102_ | _02101_;
  assign _02104_ = sel_oi_one_hot_i[106] & i[174];
  assign _02105_ = sel_oi_one_hot_i[107] & i[190];
  assign _02106_ = _02105_ | _02104_;
  assign _02107_ = _02106_ | _02103_;
  assign _02108_ = sel_oi_one_hot_i[108] & i[206];
  assign _02109_ = sel_oi_one_hot_i[109] & i[222];
  assign _02110_ = _02109_ | _02108_;
  assign _02111_ = sel_oi_one_hot_i[110] & i[238];
  assign _02112_ = sel_oi_one_hot_i[111] & i[254];
  assign _02113_ = _02112_ | _02111_;
  assign _02114_ = _02113_ | _02110_;
  assign _02115_ = _02114_ | _02107_;
  assign o[110] = _02115_ | _02100_;
  assign _02116_ = sel_oi_one_hot_i[96] & i[13];
  assign _02117_ = sel_oi_one_hot_i[97] & i[29];
  assign _02118_ = _02117_ | _02116_;
  assign _02119_ = sel_oi_one_hot_i[98] & i[45];
  assign _02120_ = sel_oi_one_hot_i[99] & i[61];
  assign _02121_ = _02120_ | _02119_;
  assign _02122_ = _02121_ | _02118_;
  assign _02123_ = sel_oi_one_hot_i[100] & i[77];
  assign _02124_ = sel_oi_one_hot_i[101] & i[93];
  assign _02125_ = _02124_ | _02123_;
  assign _02126_ = sel_oi_one_hot_i[102] & i[109];
  assign _02127_ = sel_oi_one_hot_i[103] & i[125];
  assign _02128_ = _02127_ | _02126_;
  assign _02129_ = _02128_ | _02125_;
  assign _02130_ = _02129_ | _02122_;
  assign _02131_ = sel_oi_one_hot_i[104] & i[141];
  assign _02132_ = sel_oi_one_hot_i[105] & i[157];
  assign _02133_ = _02132_ | _02131_;
  assign _02134_ = sel_oi_one_hot_i[106] & i[173];
  assign _02135_ = sel_oi_one_hot_i[107] & i[189];
  assign _02136_ = _02135_ | _02134_;
  assign _02137_ = _02136_ | _02133_;
  assign _02138_ = sel_oi_one_hot_i[108] & i[205];
  assign _02139_ = sel_oi_one_hot_i[109] & i[221];
  assign _02140_ = _02139_ | _02138_;
  assign _02141_ = sel_oi_one_hot_i[110] & i[237];
  assign _02142_ = sel_oi_one_hot_i[111] & i[253];
  assign _02143_ = _02142_ | _02141_;
  assign _02144_ = _02143_ | _02140_;
  assign _02145_ = _02144_ | _02137_;
  assign o[109] = _02145_ | _02130_;
  assign _02146_ = sel_oi_one_hot_i[96] & i[12];
  assign _02147_ = sel_oi_one_hot_i[97] & i[28];
  assign _02148_ = _02147_ | _02146_;
  assign _02149_ = sel_oi_one_hot_i[98] & i[44];
  assign _02150_ = sel_oi_one_hot_i[99] & i[60];
  assign _02151_ = _02150_ | _02149_;
  assign _02152_ = _02151_ | _02148_;
  assign _02153_ = sel_oi_one_hot_i[100] & i[76];
  assign _02154_ = sel_oi_one_hot_i[101] & i[92];
  assign _02155_ = _02154_ | _02153_;
  assign _02156_ = sel_oi_one_hot_i[102] & i[108];
  assign _02157_ = sel_oi_one_hot_i[103] & i[124];
  assign _02158_ = _02157_ | _02156_;
  assign _02159_ = _02158_ | _02155_;
  assign _02160_ = _02159_ | _02152_;
  assign _02161_ = sel_oi_one_hot_i[104] & i[140];
  assign _02162_ = sel_oi_one_hot_i[105] & i[156];
  assign _02163_ = _02162_ | _02161_;
  assign _02164_ = sel_oi_one_hot_i[106] & i[172];
  assign _02165_ = sel_oi_one_hot_i[107] & i[188];
  assign _02166_ = _02165_ | _02164_;
  assign _02167_ = _02166_ | _02163_;
  assign _02168_ = sel_oi_one_hot_i[108] & i[204];
  assign _02169_ = sel_oi_one_hot_i[109] & i[220];
  assign _02170_ = _02169_ | _02168_;
  assign _02171_ = sel_oi_one_hot_i[110] & i[236];
  assign _02172_ = sel_oi_one_hot_i[111] & i[252];
  assign _02173_ = _02172_ | _02171_;
  assign _02174_ = _02173_ | _02170_;
  assign _02175_ = _02174_ | _02167_;
  assign o[108] = _02175_ | _02160_;
  assign _02176_ = sel_oi_one_hot_i[0] & i[3];
  assign _02177_ = sel_oi_one_hot_i[1] & i[19];
  assign _02178_ = _02177_ | _02176_;
  assign _02179_ = sel_oi_one_hot_i[2] & i[35];
  assign _02180_ = sel_oi_one_hot_i[3] & i[51];
  assign _02181_ = _02180_ | _02179_;
  assign _02182_ = _02181_ | _02178_;
  assign _02183_ = sel_oi_one_hot_i[4] & i[67];
  assign _02184_ = sel_oi_one_hot_i[5] & i[83];
  assign _02185_ = _02184_ | _02183_;
  assign _02186_ = sel_oi_one_hot_i[6] & i[99];
  assign _02187_ = sel_oi_one_hot_i[7] & i[115];
  assign _02188_ = _02187_ | _02186_;
  assign _02189_ = _02188_ | _02185_;
  assign _02190_ = _02189_ | _02182_;
  assign _02191_ = sel_oi_one_hot_i[8] & i[131];
  assign _02192_ = sel_oi_one_hot_i[9] & i[147];
  assign _02193_ = _02192_ | _02191_;
  assign _02194_ = sel_oi_one_hot_i[10] & i[163];
  assign _02195_ = sel_oi_one_hot_i[11] & i[179];
  assign _02196_ = _02195_ | _02194_;
  assign _02197_ = _02196_ | _02193_;
  assign _02198_ = sel_oi_one_hot_i[12] & i[195];
  assign _02199_ = sel_oi_one_hot_i[13] & i[211];
  assign _02200_ = _02199_ | _02198_;
  assign _02201_ = sel_oi_one_hot_i[14] & i[227];
  assign _02202_ = sel_oi_one_hot_i[15] & i[243];
  assign _02203_ = _02202_ | _02201_;
  assign _02204_ = _02203_ | _02200_;
  assign _02205_ = _02204_ | _02197_;
  assign o[3] = _02205_ | _02190_;
  assign _02206_ = sel_oi_one_hot_i[96] & i[11];
  assign _02207_ = sel_oi_one_hot_i[97] & i[27];
  assign _02208_ = _02207_ | _02206_;
  assign _02209_ = sel_oi_one_hot_i[98] & i[43];
  assign _02210_ = sel_oi_one_hot_i[99] & i[59];
  assign _02211_ = _02210_ | _02209_;
  assign _02212_ = _02211_ | _02208_;
  assign _02213_ = sel_oi_one_hot_i[100] & i[75];
  assign _02214_ = sel_oi_one_hot_i[101] & i[91];
  assign _02215_ = _02214_ | _02213_;
  assign _02216_ = sel_oi_one_hot_i[102] & i[107];
  assign _02217_ = sel_oi_one_hot_i[103] & i[123];
  assign _02218_ = _02217_ | _02216_;
  assign _02219_ = _02218_ | _02215_;
  assign _02220_ = _02219_ | _02212_;
  assign _02221_ = sel_oi_one_hot_i[104] & i[139];
  assign _02222_ = sel_oi_one_hot_i[105] & i[155];
  assign _02223_ = _02222_ | _02221_;
  assign _02224_ = sel_oi_one_hot_i[106] & i[171];
  assign _02225_ = sel_oi_one_hot_i[107] & i[187];
  assign _02226_ = _02225_ | _02224_;
  assign _02227_ = _02226_ | _02223_;
  assign _02228_ = sel_oi_one_hot_i[108] & i[203];
  assign _02229_ = sel_oi_one_hot_i[109] & i[219];
  assign _02230_ = _02229_ | _02228_;
  assign _02231_ = sel_oi_one_hot_i[110] & i[235];
  assign _02232_ = sel_oi_one_hot_i[111] & i[251];
  assign _02233_ = _02232_ | _02231_;
  assign _02234_ = _02233_ | _02230_;
  assign _02235_ = _02234_ | _02227_;
  assign o[107] = _02235_ | _02220_;
  assign _02236_ = sel_oi_one_hot_i[96] & i[10];
  assign _02237_ = sel_oi_one_hot_i[97] & i[26];
  assign _02238_ = _02237_ | _02236_;
  assign _02239_ = sel_oi_one_hot_i[98] & i[42];
  assign _02240_ = sel_oi_one_hot_i[99] & i[58];
  assign _02241_ = _02240_ | _02239_;
  assign _02242_ = _02241_ | _02238_;
  assign _02243_ = sel_oi_one_hot_i[100] & i[74];
  assign _02244_ = sel_oi_one_hot_i[101] & i[90];
  assign _02245_ = _02244_ | _02243_;
  assign _02246_ = sel_oi_one_hot_i[102] & i[106];
  assign _02247_ = sel_oi_one_hot_i[103] & i[122];
  assign _02248_ = _02247_ | _02246_;
  assign _02249_ = _02248_ | _02245_;
  assign _02250_ = _02249_ | _02242_;
  assign _02251_ = sel_oi_one_hot_i[104] & i[138];
  assign _02252_ = sel_oi_one_hot_i[105] & i[154];
  assign _02253_ = _02252_ | _02251_;
  assign _02254_ = sel_oi_one_hot_i[106] & i[170];
  assign _02255_ = sel_oi_one_hot_i[107] & i[186];
  assign _02256_ = _02255_ | _02254_;
  assign _02257_ = _02256_ | _02253_;
  assign _02258_ = sel_oi_one_hot_i[108] & i[202];
  assign _02259_ = sel_oi_one_hot_i[109] & i[218];
  assign _02260_ = _02259_ | _02258_;
  assign _02261_ = sel_oi_one_hot_i[110] & i[234];
  assign _02262_ = sel_oi_one_hot_i[111] & i[250];
  assign _02263_ = _02262_ | _02261_;
  assign _02264_ = _02263_ | _02260_;
  assign _02265_ = _02264_ | _02257_;
  assign o[106] = _02265_ | _02250_;
  assign _02266_ = sel_oi_one_hot_i[96] & i[9];
  assign _02267_ = sel_oi_one_hot_i[97] & i[25];
  assign _02268_ = _02267_ | _02266_;
  assign _02269_ = sel_oi_one_hot_i[98] & i[41];
  assign _02270_ = sel_oi_one_hot_i[99] & i[57];
  assign _02271_ = _02270_ | _02269_;
  assign _02272_ = _02271_ | _02268_;
  assign _02273_ = sel_oi_one_hot_i[100] & i[73];
  assign _02274_ = sel_oi_one_hot_i[101] & i[89];
  assign _02275_ = _02274_ | _02273_;
  assign _02276_ = sel_oi_one_hot_i[102] & i[105];
  assign _02277_ = sel_oi_one_hot_i[103] & i[121];
  assign _02278_ = _02277_ | _02276_;
  assign _02279_ = _02278_ | _02275_;
  assign _02280_ = _02279_ | _02272_;
  assign _02281_ = sel_oi_one_hot_i[104] & i[137];
  assign _02282_ = sel_oi_one_hot_i[105] & i[153];
  assign _02283_ = _02282_ | _02281_;
  assign _02284_ = sel_oi_one_hot_i[106] & i[169];
  assign _02285_ = sel_oi_one_hot_i[107] & i[185];
  assign _02286_ = _02285_ | _02284_;
  assign _02287_ = _02286_ | _02283_;
  assign _02288_ = sel_oi_one_hot_i[108] & i[201];
  assign _02289_ = sel_oi_one_hot_i[109] & i[217];
  assign _02290_ = _02289_ | _02288_;
  assign _02291_ = sel_oi_one_hot_i[110] & i[233];
  assign _02292_ = sel_oi_one_hot_i[111] & i[249];
  assign _02293_ = _02292_ | _02291_;
  assign _02294_ = _02293_ | _02290_;
  assign _02295_ = _02294_ | _02287_;
  assign o[105] = _02295_ | _02280_;
  assign _02296_ = sel_oi_one_hot_i[96] & i[8];
  assign _02297_ = sel_oi_one_hot_i[97] & i[24];
  assign _02298_ = _02297_ | _02296_;
  assign _02299_ = sel_oi_one_hot_i[98] & i[40];
  assign _02300_ = sel_oi_one_hot_i[99] & i[56];
  assign _02301_ = _02300_ | _02299_;
  assign _02302_ = _02301_ | _02298_;
  assign _02303_ = sel_oi_one_hot_i[100] & i[72];
  assign _02304_ = sel_oi_one_hot_i[101] & i[88];
  assign _02305_ = _02304_ | _02303_;
  assign _02306_ = sel_oi_one_hot_i[102] & i[104];
  assign _02307_ = sel_oi_one_hot_i[103] & i[120];
  assign _02308_ = _02307_ | _02306_;
  assign _02309_ = _02308_ | _02305_;
  assign _02310_ = _02309_ | _02302_;
  assign _02311_ = sel_oi_one_hot_i[104] & i[136];
  assign _02312_ = sel_oi_one_hot_i[105] & i[152];
  assign _02313_ = _02312_ | _02311_;
  assign _02314_ = sel_oi_one_hot_i[106] & i[168];
  assign _02315_ = sel_oi_one_hot_i[107] & i[184];
  assign _02316_ = _02315_ | _02314_;
  assign _02317_ = _02316_ | _02313_;
  assign _02318_ = sel_oi_one_hot_i[108] & i[200];
  assign _02319_ = sel_oi_one_hot_i[109] & i[216];
  assign _02320_ = _02319_ | _02318_;
  assign _02321_ = sel_oi_one_hot_i[110] & i[232];
  assign _02322_ = sel_oi_one_hot_i[111] & i[248];
  assign _02323_ = _02322_ | _02321_;
  assign _02324_ = _02323_ | _02320_;
  assign _02325_ = _02324_ | _02317_;
  assign o[104] = _02325_ | _02310_;
  assign _02326_ = sel_oi_one_hot_i[96] & i[7];
  assign _02327_ = sel_oi_one_hot_i[97] & i[23];
  assign _02328_ = _02327_ | _02326_;
  assign _02329_ = sel_oi_one_hot_i[98] & i[39];
  assign _02330_ = sel_oi_one_hot_i[99] & i[55];
  assign _02331_ = _02330_ | _02329_;
  assign _02332_ = _02331_ | _02328_;
  assign _02333_ = sel_oi_one_hot_i[100] & i[71];
  assign _02334_ = sel_oi_one_hot_i[101] & i[87];
  assign _02335_ = _02334_ | _02333_;
  assign _02336_ = sel_oi_one_hot_i[102] & i[103];
  assign _02337_ = sel_oi_one_hot_i[103] & i[119];
  assign _02338_ = _02337_ | _02336_;
  assign _02339_ = _02338_ | _02335_;
  assign _02340_ = _02339_ | _02332_;
  assign _02341_ = sel_oi_one_hot_i[104] & i[135];
  assign _02342_ = sel_oi_one_hot_i[105] & i[151];
  assign _02343_ = _02342_ | _02341_;
  assign _02344_ = sel_oi_one_hot_i[106] & i[167];
  assign _02345_ = sel_oi_one_hot_i[107] & i[183];
  assign _02346_ = _02345_ | _02344_;
  assign _02347_ = _02346_ | _02343_;
  assign _02348_ = sel_oi_one_hot_i[108] & i[199];
  assign _02349_ = sel_oi_one_hot_i[109] & i[215];
  assign _02350_ = _02349_ | _02348_;
  assign _02351_ = sel_oi_one_hot_i[110] & i[231];
  assign _02352_ = sel_oi_one_hot_i[111] & i[247];
  assign _02353_ = _02352_ | _02351_;
  assign _02354_ = _02353_ | _02350_;
  assign _02355_ = _02354_ | _02347_;
  assign o[103] = _02355_ | _02340_;
  assign _02356_ = sel_oi_one_hot_i[96] & i[6];
  assign _02357_ = sel_oi_one_hot_i[97] & i[22];
  assign _02358_ = _02357_ | _02356_;
  assign _02359_ = sel_oi_one_hot_i[98] & i[38];
  assign _02360_ = sel_oi_one_hot_i[99] & i[54];
  assign _02361_ = _02360_ | _02359_;
  assign _02362_ = _02361_ | _02358_;
  assign _02363_ = sel_oi_one_hot_i[100] & i[70];
  assign _02364_ = sel_oi_one_hot_i[101] & i[86];
  assign _02365_ = _02364_ | _02363_;
  assign _02366_ = sel_oi_one_hot_i[102] & i[102];
  assign _02367_ = sel_oi_one_hot_i[103] & i[118];
  assign _02368_ = _02367_ | _02366_;
  assign _02369_ = _02368_ | _02365_;
  assign _02370_ = _02369_ | _02362_;
  assign _02371_ = sel_oi_one_hot_i[104] & i[134];
  assign _02372_ = sel_oi_one_hot_i[105] & i[150];
  assign _02373_ = _02372_ | _02371_;
  assign _02374_ = sel_oi_one_hot_i[106] & i[166];
  assign _02375_ = sel_oi_one_hot_i[107] & i[182];
  assign _02376_ = _02375_ | _02374_;
  assign _02377_ = _02376_ | _02373_;
  assign _02378_ = sel_oi_one_hot_i[108] & i[198];
  assign _02379_ = sel_oi_one_hot_i[109] & i[214];
  assign _02380_ = _02379_ | _02378_;
  assign _02381_ = sel_oi_one_hot_i[110] & i[230];
  assign _02382_ = sel_oi_one_hot_i[111] & i[246];
  assign _02383_ = _02382_ | _02381_;
  assign _02384_ = _02383_ | _02380_;
  assign _02385_ = _02384_ | _02377_;
  assign o[102] = _02385_ | _02370_;
  assign _02386_ = sel_oi_one_hot_i[96] & i[5];
  assign _02387_ = sel_oi_one_hot_i[97] & i[21];
  assign _02388_ = _02387_ | _02386_;
  assign _02389_ = sel_oi_one_hot_i[98] & i[37];
  assign _02390_ = sel_oi_one_hot_i[99] & i[53];
  assign _02391_ = _02390_ | _02389_;
  assign _02392_ = _02391_ | _02388_;
  assign _02393_ = sel_oi_one_hot_i[100] & i[69];
  assign _02394_ = sel_oi_one_hot_i[101] & i[85];
  assign _02395_ = _02394_ | _02393_;
  assign _02396_ = sel_oi_one_hot_i[102] & i[101];
  assign _02397_ = sel_oi_one_hot_i[103] & i[117];
  assign _02398_ = _02397_ | _02396_;
  assign _02399_ = _02398_ | _02395_;
  assign _02400_ = _02399_ | _02392_;
  assign _02401_ = sel_oi_one_hot_i[104] & i[133];
  assign _02402_ = sel_oi_one_hot_i[105] & i[149];
  assign _02403_ = _02402_ | _02401_;
  assign _02404_ = sel_oi_one_hot_i[106] & i[165];
  assign _02405_ = sel_oi_one_hot_i[107] & i[181];
  assign _02406_ = _02405_ | _02404_;
  assign _02407_ = _02406_ | _02403_;
  assign _02408_ = sel_oi_one_hot_i[108] & i[197];
  assign _02409_ = sel_oi_one_hot_i[109] & i[213];
  assign _02410_ = _02409_ | _02408_;
  assign _02411_ = sel_oi_one_hot_i[110] & i[229];
  assign _02412_ = sel_oi_one_hot_i[111] & i[245];
  assign _02413_ = _02412_ | _02411_;
  assign _02414_ = _02413_ | _02410_;
  assign _02415_ = _02414_ | _02407_;
  assign o[101] = _02415_ | _02400_;
  assign _02416_ = sel_oi_one_hot_i[96] & i[4];
  assign _02417_ = sel_oi_one_hot_i[97] & i[20];
  assign _02418_ = _02417_ | _02416_;
  assign _02419_ = sel_oi_one_hot_i[98] & i[36];
  assign _02420_ = sel_oi_one_hot_i[99] & i[52];
  assign _02421_ = _02420_ | _02419_;
  assign _02422_ = _02421_ | _02418_;
  assign _02423_ = sel_oi_one_hot_i[100] & i[68];
  assign _02424_ = sel_oi_one_hot_i[101] & i[84];
  assign _02425_ = _02424_ | _02423_;
  assign _02426_ = sel_oi_one_hot_i[102] & i[100];
  assign _02427_ = sel_oi_one_hot_i[103] & i[116];
  assign _02428_ = _02427_ | _02426_;
  assign _02429_ = _02428_ | _02425_;
  assign _02430_ = _02429_ | _02422_;
  assign _02431_ = sel_oi_one_hot_i[104] & i[132];
  assign _02432_ = sel_oi_one_hot_i[105] & i[148];
  assign _02433_ = _02432_ | _02431_;
  assign _02434_ = sel_oi_one_hot_i[106] & i[164];
  assign _02435_ = sel_oi_one_hot_i[107] & i[180];
  assign _02436_ = _02435_ | _02434_;
  assign _02437_ = _02436_ | _02433_;
  assign _02438_ = sel_oi_one_hot_i[108] & i[196];
  assign _02439_ = sel_oi_one_hot_i[109] & i[212];
  assign _02440_ = _02439_ | _02438_;
  assign _02441_ = sel_oi_one_hot_i[110] & i[228];
  assign _02442_ = sel_oi_one_hot_i[111] & i[244];
  assign _02443_ = _02442_ | _02441_;
  assign _02444_ = _02443_ | _02440_;
  assign _02445_ = _02444_ | _02437_;
  assign o[100] = _02445_ | _02430_;
  assign _02446_ = sel_oi_one_hot_i[96] & i[3];
  assign _02447_ = sel_oi_one_hot_i[97] & i[19];
  assign _02448_ = _02447_ | _02446_;
  assign _02449_ = sel_oi_one_hot_i[98] & i[35];
  assign _02450_ = sel_oi_one_hot_i[99] & i[51];
  assign _02451_ = _02450_ | _02449_;
  assign _02452_ = _02451_ | _02448_;
  assign _02453_ = sel_oi_one_hot_i[100] & i[67];
  assign _02454_ = sel_oi_one_hot_i[101] & i[83];
  assign _02455_ = _02454_ | _02453_;
  assign _02456_ = sel_oi_one_hot_i[102] & i[99];
  assign _02457_ = sel_oi_one_hot_i[103] & i[115];
  assign _02458_ = _02457_ | _02456_;
  assign _02459_ = _02458_ | _02455_;
  assign _02460_ = _02459_ | _02452_;
  assign _02461_ = sel_oi_one_hot_i[104] & i[131];
  assign _02462_ = sel_oi_one_hot_i[105] & i[147];
  assign _02463_ = _02462_ | _02461_;
  assign _02464_ = sel_oi_one_hot_i[106] & i[163];
  assign _02465_ = sel_oi_one_hot_i[107] & i[179];
  assign _02466_ = _02465_ | _02464_;
  assign _02467_ = _02466_ | _02463_;
  assign _02468_ = sel_oi_one_hot_i[108] & i[195];
  assign _02469_ = sel_oi_one_hot_i[109] & i[211];
  assign _02470_ = _02469_ | _02468_;
  assign _02471_ = sel_oi_one_hot_i[110] & i[227];
  assign _02472_ = sel_oi_one_hot_i[111] & i[243];
  assign _02473_ = _02472_ | _02471_;
  assign _02474_ = _02473_ | _02470_;
  assign _02475_ = _02474_ | _02467_;
  assign o[99] = _02475_ | _02460_;
  assign _02476_ = sel_oi_one_hot_i[96] & i[2];
  assign _02477_ = sel_oi_one_hot_i[97] & i[18];
  assign _02478_ = _02477_ | _02476_;
  assign _02479_ = sel_oi_one_hot_i[98] & i[34];
  assign _02480_ = sel_oi_one_hot_i[99] & i[50];
  assign _02481_ = _02480_ | _02479_;
  assign _02482_ = _02481_ | _02478_;
  assign _02483_ = sel_oi_one_hot_i[100] & i[66];
  assign _02484_ = sel_oi_one_hot_i[101] & i[82];
  assign _02485_ = _02484_ | _02483_;
  assign _02486_ = sel_oi_one_hot_i[102] & i[98];
  assign _02487_ = sel_oi_one_hot_i[103] & i[114];
  assign _02488_ = _02487_ | _02486_;
  assign _02489_ = _02488_ | _02485_;
  assign _02490_ = _02489_ | _02482_;
  assign _02491_ = sel_oi_one_hot_i[104] & i[130];
  assign _02492_ = sel_oi_one_hot_i[105] & i[146];
  assign _02493_ = _02492_ | _02491_;
  assign _02494_ = sel_oi_one_hot_i[106] & i[162];
  assign _02495_ = sel_oi_one_hot_i[107] & i[178];
  assign _02496_ = _02495_ | _02494_;
  assign _02497_ = _02496_ | _02493_;
  assign _02498_ = sel_oi_one_hot_i[108] & i[194];
  assign _02499_ = sel_oi_one_hot_i[109] & i[210];
  assign _02500_ = _02499_ | _02498_;
  assign _02501_ = sel_oi_one_hot_i[110] & i[226];
  assign _02502_ = sel_oi_one_hot_i[111] & i[242];
  assign _02503_ = _02502_ | _02501_;
  assign _02504_ = _02503_ | _02500_;
  assign _02505_ = _02504_ | _02497_;
  assign o[98] = _02505_ | _02490_;
  assign _02506_ = sel_oi_one_hot_i[0] & i[2];
  assign _02507_ = sel_oi_one_hot_i[1] & i[18];
  assign _02508_ = _02507_ | _02506_;
  assign _02509_ = sel_oi_one_hot_i[2] & i[34];
  assign _02510_ = sel_oi_one_hot_i[3] & i[50];
  assign _02511_ = _02510_ | _02509_;
  assign _02512_ = _02511_ | _02508_;
  assign _02513_ = sel_oi_one_hot_i[4] & i[66];
  assign _02514_ = sel_oi_one_hot_i[5] & i[82];
  assign _02515_ = _02514_ | _02513_;
  assign _02516_ = sel_oi_one_hot_i[6] & i[98];
  assign _02517_ = sel_oi_one_hot_i[7] & i[114];
  assign _02518_ = _02517_ | _02516_;
  assign _02519_ = _02518_ | _02515_;
  assign _02520_ = _02519_ | _02512_;
  assign _02521_ = sel_oi_one_hot_i[8] & i[130];
  assign _02522_ = sel_oi_one_hot_i[9] & i[146];
  assign _02523_ = _02522_ | _02521_;
  assign _02524_ = sel_oi_one_hot_i[10] & i[162];
  assign _02525_ = sel_oi_one_hot_i[11] & i[178];
  assign _02526_ = _02525_ | _02524_;
  assign _02527_ = _02526_ | _02523_;
  assign _02528_ = sel_oi_one_hot_i[12] & i[194];
  assign _02529_ = sel_oi_one_hot_i[13] & i[210];
  assign _02530_ = _02529_ | _02528_;
  assign _02531_ = sel_oi_one_hot_i[14] & i[226];
  assign _02532_ = sel_oi_one_hot_i[15] & i[242];
  assign _02533_ = _02532_ | _02531_;
  assign _02534_ = _02533_ | _02530_;
  assign _02535_ = _02534_ | _02527_;
  assign o[2] = _02535_ | _02520_;
  assign _02536_ = sel_oi_one_hot_i[96] & i[1];
  assign _02537_ = sel_oi_one_hot_i[97] & i[17];
  assign _02538_ = _02537_ | _02536_;
  assign _02539_ = sel_oi_one_hot_i[98] & i[33];
  assign _02540_ = sel_oi_one_hot_i[99] & i[49];
  assign _02541_ = _02540_ | _02539_;
  assign _02542_ = _02541_ | _02538_;
  assign _02543_ = sel_oi_one_hot_i[100] & i[65];
  assign _02544_ = sel_oi_one_hot_i[101] & i[81];
  assign _02545_ = _02544_ | _02543_;
  assign _02546_ = sel_oi_one_hot_i[102] & i[97];
  assign _02547_ = sel_oi_one_hot_i[103] & i[113];
  assign _02548_ = _02547_ | _02546_;
  assign _02549_ = _02548_ | _02545_;
  assign _02550_ = _02549_ | _02542_;
  assign _02551_ = sel_oi_one_hot_i[104] & i[129];
  assign _02552_ = sel_oi_one_hot_i[105] & i[145];
  assign _02553_ = _02552_ | _02551_;
  assign _02554_ = sel_oi_one_hot_i[106] & i[161];
  assign _02555_ = sel_oi_one_hot_i[107] & i[177];
  assign _02556_ = _02555_ | _02554_;
  assign _02557_ = _02556_ | _02553_;
  assign _02558_ = sel_oi_one_hot_i[108] & i[193];
  assign _02559_ = sel_oi_one_hot_i[109] & i[209];
  assign _02560_ = _02559_ | _02558_;
  assign _02561_ = sel_oi_one_hot_i[110] & i[225];
  assign _02562_ = sel_oi_one_hot_i[111] & i[241];
  assign _02563_ = _02562_ | _02561_;
  assign _02564_ = _02563_ | _02560_;
  assign _02565_ = _02564_ | _02557_;
  assign o[97] = _02565_ | _02550_;
  assign _02566_ = sel_oi_one_hot_i[96] & i[0];
  assign _02567_ = sel_oi_one_hot_i[97] & i[16];
  assign _02568_ = _02567_ | _02566_;
  assign _02569_ = sel_oi_one_hot_i[98] & i[32];
  assign _02570_ = sel_oi_one_hot_i[99] & i[48];
  assign _02571_ = _02570_ | _02569_;
  assign _02572_ = _02571_ | _02568_;
  assign _02573_ = sel_oi_one_hot_i[100] & i[64];
  assign _02574_ = sel_oi_one_hot_i[101] & i[80];
  assign _02575_ = _02574_ | _02573_;
  assign _02576_ = sel_oi_one_hot_i[102] & i[96];
  assign _02577_ = sel_oi_one_hot_i[103] & i[112];
  assign _02578_ = _02577_ | _02576_;
  assign _02579_ = _02578_ | _02575_;
  assign _02580_ = _02579_ | _02572_;
  assign _02581_ = sel_oi_one_hot_i[104] & i[128];
  assign _02582_ = sel_oi_one_hot_i[105] & i[144];
  assign _02583_ = _02582_ | _02581_;
  assign _02584_ = sel_oi_one_hot_i[106] & i[160];
  assign _02585_ = sel_oi_one_hot_i[107] & i[176];
  assign _02586_ = _02585_ | _02584_;
  assign _02587_ = _02586_ | _02583_;
  assign _02588_ = sel_oi_one_hot_i[108] & i[192];
  assign _02589_ = sel_oi_one_hot_i[109] & i[208];
  assign _02590_ = _02589_ | _02588_;
  assign _02591_ = sel_oi_one_hot_i[110] & i[224];
  assign _02592_ = sel_oi_one_hot_i[111] & i[240];
  assign _02593_ = _02592_ | _02591_;
  assign _02594_ = _02593_ | _02590_;
  assign _02595_ = _02594_ | _02587_;
  assign o[96] = _02595_ | _02580_;
  assign _02596_ = sel_oi_one_hot_i[0] & i[1];
  assign _02597_ = sel_oi_one_hot_i[1] & i[17];
  assign _02598_ = _02597_ | _02596_;
  assign _02599_ = sel_oi_one_hot_i[2] & i[33];
  assign _02600_ = sel_oi_one_hot_i[3] & i[49];
  assign _02601_ = _02600_ | _02599_;
  assign _02602_ = _02601_ | _02598_;
  assign _02603_ = sel_oi_one_hot_i[4] & i[65];
  assign _02604_ = sel_oi_one_hot_i[5] & i[81];
  assign _02605_ = _02604_ | _02603_;
  assign _02606_ = sel_oi_one_hot_i[6] & i[97];
  assign _02607_ = sel_oi_one_hot_i[7] & i[113];
  assign _02608_ = _02607_ | _02606_;
  assign _02609_ = _02608_ | _02605_;
  assign _02610_ = _02609_ | _02602_;
  assign _02611_ = sel_oi_one_hot_i[8] & i[129];
  assign _02612_ = sel_oi_one_hot_i[9] & i[145];
  assign _02613_ = _02612_ | _02611_;
  assign _02614_ = sel_oi_one_hot_i[10] & i[161];
  assign _02615_ = sel_oi_one_hot_i[11] & i[177];
  assign _02616_ = _02615_ | _02614_;
  assign _02617_ = _02616_ | _02613_;
  assign _02618_ = sel_oi_one_hot_i[12] & i[193];
  assign _02619_ = sel_oi_one_hot_i[13] & i[209];
  assign _02620_ = _02619_ | _02618_;
  assign _02621_ = sel_oi_one_hot_i[14] & i[225];
  assign _02622_ = sel_oi_one_hot_i[15] & i[241];
  assign _02623_ = _02622_ | _02621_;
  assign _02624_ = _02623_ | _02620_;
  assign _02625_ = _02624_ | _02617_;
  assign o[1] = _02625_ | _02610_;
  assign _02626_ = sel_oi_one_hot_i[112] & i[15];
  assign _02627_ = sel_oi_one_hot_i[113] & i[31];
  assign _02628_ = _02627_ | _02626_;
  assign _02629_ = sel_oi_one_hot_i[114] & i[47];
  assign _02630_ = sel_oi_one_hot_i[115] & i[63];
  assign _02631_ = _02630_ | _02629_;
  assign _02632_ = _02631_ | _02628_;
  assign _02633_ = sel_oi_one_hot_i[116] & i[79];
  assign _02634_ = sel_oi_one_hot_i[117] & i[95];
  assign _02635_ = _02634_ | _02633_;
  assign _02636_ = sel_oi_one_hot_i[118] & i[111];
  assign _02637_ = sel_oi_one_hot_i[119] & i[127];
  assign _02638_ = _02637_ | _02636_;
  assign _02639_ = _02638_ | _02635_;
  assign _02640_ = _02639_ | _02632_;
  assign _02641_ = sel_oi_one_hot_i[120] & i[143];
  assign _02642_ = sel_oi_one_hot_i[121] & i[159];
  assign _02643_ = _02642_ | _02641_;
  assign _02644_ = sel_oi_one_hot_i[122] & i[175];
  assign _02645_ = sel_oi_one_hot_i[123] & i[191];
  assign _02646_ = _02645_ | _02644_;
  assign _02647_ = _02646_ | _02643_;
  assign _02648_ = sel_oi_one_hot_i[124] & i[207];
  assign _02649_ = sel_oi_one_hot_i[125] & i[223];
  assign _02650_ = _02649_ | _02648_;
  assign _02651_ = sel_oi_one_hot_i[126] & i[239];
  assign _02652_ = sel_oi_one_hot_i[127] & i[255];
  assign _02653_ = _02652_ | _02651_;
  assign _02654_ = _02653_ | _02650_;
  assign _02655_ = _02654_ | _02647_;
  assign o[127] = _02655_ | _02640_;
  assign _02656_ = sel_oi_one_hot_i[112] & i[14];
  assign _02657_ = sel_oi_one_hot_i[113] & i[30];
  assign _02658_ = _02657_ | _02656_;
  assign _02659_ = sel_oi_one_hot_i[114] & i[46];
  assign _02660_ = sel_oi_one_hot_i[115] & i[62];
  assign _02661_ = _02660_ | _02659_;
  assign _02662_ = _02661_ | _02658_;
  assign _02663_ = sel_oi_one_hot_i[116] & i[78];
  assign _02664_ = sel_oi_one_hot_i[117] & i[94];
  assign _02665_ = _02664_ | _02663_;
  assign _02666_ = sel_oi_one_hot_i[118] & i[110];
  assign _02667_ = sel_oi_one_hot_i[119] & i[126];
  assign _02668_ = _02667_ | _02666_;
  assign _02669_ = _02668_ | _02665_;
  assign _02670_ = _02669_ | _02662_;
  assign _02671_ = sel_oi_one_hot_i[120] & i[142];
  assign _02672_ = sel_oi_one_hot_i[121] & i[158];
  assign _02673_ = _02672_ | _02671_;
  assign _02674_ = sel_oi_one_hot_i[122] & i[174];
  assign _02675_ = sel_oi_one_hot_i[123] & i[190];
  assign _02676_ = _02675_ | _02674_;
  assign _02677_ = _02676_ | _02673_;
  assign _02678_ = sel_oi_one_hot_i[124] & i[206];
  assign _02679_ = sel_oi_one_hot_i[125] & i[222];
  assign _02680_ = _02679_ | _02678_;
  assign _02681_ = sel_oi_one_hot_i[126] & i[238];
  assign _02682_ = sel_oi_one_hot_i[127] & i[254];
  assign _02683_ = _02682_ | _02681_;
  assign _02684_ = _02683_ | _02680_;
  assign _02685_ = _02684_ | _02677_;
  assign o[126] = _02685_ | _02670_;
  assign _02686_ = sel_oi_one_hot_i[112] & i[13];
  assign _02687_ = sel_oi_one_hot_i[113] & i[29];
  assign _02688_ = _02687_ | _02686_;
  assign _02689_ = sel_oi_one_hot_i[114] & i[45];
  assign _02690_ = sel_oi_one_hot_i[115] & i[61];
  assign _02691_ = _02690_ | _02689_;
  assign _02692_ = _02691_ | _02688_;
  assign _02693_ = sel_oi_one_hot_i[116] & i[77];
  assign _02694_ = sel_oi_one_hot_i[117] & i[93];
  assign _02695_ = _02694_ | _02693_;
  assign _02696_ = sel_oi_one_hot_i[118] & i[109];
  assign _02697_ = sel_oi_one_hot_i[119] & i[125];
  assign _02698_ = _02697_ | _02696_;
  assign _02699_ = _02698_ | _02695_;
  assign _02700_ = _02699_ | _02692_;
  assign _02701_ = sel_oi_one_hot_i[120] & i[141];
  assign _02702_ = sel_oi_one_hot_i[121] & i[157];
  assign _02703_ = _02702_ | _02701_;
  assign _02704_ = sel_oi_one_hot_i[122] & i[173];
  assign _02705_ = sel_oi_one_hot_i[123] & i[189];
  assign _02706_ = _02705_ | _02704_;
  assign _02707_ = _02706_ | _02703_;
  assign _02708_ = sel_oi_one_hot_i[124] & i[205];
  assign _02709_ = sel_oi_one_hot_i[125] & i[221];
  assign _02710_ = _02709_ | _02708_;
  assign _02711_ = sel_oi_one_hot_i[126] & i[237];
  assign _02712_ = sel_oi_one_hot_i[127] & i[253];
  assign _02713_ = _02712_ | _02711_;
  assign _02714_ = _02713_ | _02710_;
  assign _02715_ = _02714_ | _02707_;
  assign o[125] = _02715_ | _02700_;
  assign _02716_ = sel_oi_one_hot_i[112] & i[12];
  assign _02717_ = sel_oi_one_hot_i[113] & i[28];
  assign _02718_ = _02717_ | _02716_;
  assign _02719_ = sel_oi_one_hot_i[114] & i[44];
  assign _02720_ = sel_oi_one_hot_i[115] & i[60];
  assign _02721_ = _02720_ | _02719_;
  assign _02722_ = _02721_ | _02718_;
  assign _02723_ = sel_oi_one_hot_i[116] & i[76];
  assign _02724_ = sel_oi_one_hot_i[117] & i[92];
  assign _02725_ = _02724_ | _02723_;
  assign _02726_ = sel_oi_one_hot_i[118] & i[108];
  assign _02727_ = sel_oi_one_hot_i[119] & i[124];
  assign _02728_ = _02727_ | _02726_;
  assign _02729_ = _02728_ | _02725_;
  assign _02730_ = _02729_ | _02722_;
  assign _02731_ = sel_oi_one_hot_i[120] & i[140];
  assign _02732_ = sel_oi_one_hot_i[121] & i[156];
  assign _02733_ = _02732_ | _02731_;
  assign _02734_ = sel_oi_one_hot_i[122] & i[172];
  assign _02735_ = sel_oi_one_hot_i[123] & i[188];
  assign _02736_ = _02735_ | _02734_;
  assign _02737_ = _02736_ | _02733_;
  assign _02738_ = sel_oi_one_hot_i[124] & i[204];
  assign _02739_ = sel_oi_one_hot_i[125] & i[220];
  assign _02740_ = _02739_ | _02738_;
  assign _02741_ = sel_oi_one_hot_i[126] & i[236];
  assign _02742_ = sel_oi_one_hot_i[127] & i[252];
  assign _02743_ = _02742_ | _02741_;
  assign _02744_ = _02743_ | _02740_;
  assign _02745_ = _02744_ | _02737_;
  assign o[124] = _02745_ | _02730_;
  assign _02746_ = sel_oi_one_hot_i[112] & i[11];
  assign _02747_ = sel_oi_one_hot_i[113] & i[27];
  assign _02748_ = _02747_ | _02746_;
  assign _02749_ = sel_oi_one_hot_i[114] & i[43];
  assign _02750_ = sel_oi_one_hot_i[115] & i[59];
  assign _02751_ = _02750_ | _02749_;
  assign _02752_ = _02751_ | _02748_;
  assign _02753_ = sel_oi_one_hot_i[116] & i[75];
  assign _02754_ = sel_oi_one_hot_i[117] & i[91];
  assign _02755_ = _02754_ | _02753_;
  assign _02756_ = sel_oi_one_hot_i[118] & i[107];
  assign _02757_ = sel_oi_one_hot_i[119] & i[123];
  assign _02758_ = _02757_ | _02756_;
  assign _02759_ = _02758_ | _02755_;
  assign _02760_ = _02759_ | _02752_;
  assign _02761_ = sel_oi_one_hot_i[120] & i[139];
  assign _02762_ = sel_oi_one_hot_i[121] & i[155];
  assign _02763_ = _02762_ | _02761_;
  assign _02764_ = sel_oi_one_hot_i[122] & i[171];
  assign _02765_ = sel_oi_one_hot_i[123] & i[187];
  assign _02766_ = _02765_ | _02764_;
  assign _02767_ = _02766_ | _02763_;
  assign _02768_ = sel_oi_one_hot_i[124] & i[203];
  assign _02769_ = sel_oi_one_hot_i[125] & i[219];
  assign _02770_ = _02769_ | _02768_;
  assign _02771_ = sel_oi_one_hot_i[126] & i[235];
  assign _02772_ = sel_oi_one_hot_i[127] & i[251];
  assign _02773_ = _02772_ | _02771_;
  assign _02774_ = _02773_ | _02770_;
  assign _02775_ = _02774_ | _02767_;
  assign o[123] = _02775_ | _02760_;
  assign _02776_ = sel_oi_one_hot_i[0] & i[0];
  assign _02777_ = sel_oi_one_hot_i[1] & i[16];
  assign _02778_ = _02777_ | _02776_;
  assign _02779_ = sel_oi_one_hot_i[2] & i[32];
  assign _02780_ = sel_oi_one_hot_i[3] & i[48];
  assign _02781_ = _02780_ | _02779_;
  assign _02782_ = _02781_ | _02778_;
  assign _02783_ = sel_oi_one_hot_i[4] & i[64];
  assign _02784_ = sel_oi_one_hot_i[5] & i[80];
  assign _02785_ = _02784_ | _02783_;
  assign _02786_ = sel_oi_one_hot_i[6] & i[96];
  assign _02787_ = sel_oi_one_hot_i[7] & i[112];
  assign _02788_ = _02787_ | _02786_;
  assign _02789_ = _02788_ | _02785_;
  assign _02790_ = _02789_ | _02782_;
  assign _02791_ = sel_oi_one_hot_i[8] & i[128];
  assign _02792_ = sel_oi_one_hot_i[9] & i[144];
  assign _02793_ = _02792_ | _02791_;
  assign _02794_ = sel_oi_one_hot_i[10] & i[160];
  assign _02795_ = sel_oi_one_hot_i[11] & i[176];
  assign _02796_ = _02795_ | _02794_;
  assign _02797_ = _02796_ | _02793_;
  assign _02798_ = sel_oi_one_hot_i[12] & i[192];
  assign _02799_ = sel_oi_one_hot_i[13] & i[208];
  assign _02800_ = _02799_ | _02798_;
  assign _02801_ = sel_oi_one_hot_i[14] & i[224];
  assign _02802_ = sel_oi_one_hot_i[15] & i[240];
  assign _02803_ = _02802_ | _02801_;
  assign _02804_ = _02803_ | _02800_;
  assign _02805_ = _02804_ | _02797_;
  assign o[0] = _02805_ | _02790_;
  assign _02806_ = sel_oi_one_hot_i[112] & i[10];
  assign _02807_ = sel_oi_one_hot_i[113] & i[26];
  assign _02808_ = _02807_ | _02806_;
  assign _02809_ = sel_oi_one_hot_i[114] & i[42];
  assign _02810_ = sel_oi_one_hot_i[115] & i[58];
  assign _02811_ = _02810_ | _02809_;
  assign _02812_ = _02811_ | _02808_;
  assign _02813_ = sel_oi_one_hot_i[116] & i[74];
  assign _02814_ = sel_oi_one_hot_i[117] & i[90];
  assign _02815_ = _02814_ | _02813_;
  assign _02816_ = sel_oi_one_hot_i[118] & i[106];
  assign _02817_ = sel_oi_one_hot_i[119] & i[122];
  assign _02818_ = _02817_ | _02816_;
  assign _02819_ = _02818_ | _02815_;
  assign _02820_ = _02819_ | _02812_;
  assign _02821_ = sel_oi_one_hot_i[120] & i[138];
  assign _02822_ = sel_oi_one_hot_i[121] & i[154];
  assign _02823_ = _02822_ | _02821_;
  assign _02824_ = sel_oi_one_hot_i[122] & i[170];
  assign _02825_ = sel_oi_one_hot_i[123] & i[186];
  assign _02826_ = _02825_ | _02824_;
  assign _02827_ = _02826_ | _02823_;
  assign _02828_ = sel_oi_one_hot_i[124] & i[202];
  assign _02829_ = sel_oi_one_hot_i[125] & i[218];
  assign _02830_ = _02829_ | _02828_;
  assign _02831_ = sel_oi_one_hot_i[126] & i[234];
  assign _02832_ = sel_oi_one_hot_i[127] & i[250];
  assign _02833_ = _02832_ | _02831_;
  assign _02834_ = _02833_ | _02830_;
  assign _02835_ = _02834_ | _02827_;
  assign o[122] = _02835_ | _02820_;
  assign _02836_ = sel_oi_one_hot_i[112] & i[9];
  assign _02837_ = sel_oi_one_hot_i[113] & i[25];
  assign _02838_ = _02837_ | _02836_;
  assign _02839_ = sel_oi_one_hot_i[114] & i[41];
  assign _02840_ = sel_oi_one_hot_i[115] & i[57];
  assign _02841_ = _02840_ | _02839_;
  assign _02842_ = _02841_ | _02838_;
  assign _02843_ = sel_oi_one_hot_i[116] & i[73];
  assign _02844_ = sel_oi_one_hot_i[117] & i[89];
  assign _02845_ = _02844_ | _02843_;
  assign _02846_ = sel_oi_one_hot_i[118] & i[105];
  assign _02847_ = sel_oi_one_hot_i[119] & i[121];
  assign _02848_ = _02847_ | _02846_;
  assign _02849_ = _02848_ | _02845_;
  assign _02850_ = _02849_ | _02842_;
  assign _02851_ = sel_oi_one_hot_i[120] & i[137];
  assign _02852_ = sel_oi_one_hot_i[121] & i[153];
  assign _02853_ = _02852_ | _02851_;
  assign _02854_ = sel_oi_one_hot_i[122] & i[169];
  assign _02855_ = sel_oi_one_hot_i[123] & i[185];
  assign _02856_ = _02855_ | _02854_;
  assign _02857_ = _02856_ | _02853_;
  assign _02858_ = sel_oi_one_hot_i[124] & i[201];
  assign _02859_ = sel_oi_one_hot_i[125] & i[217];
  assign _02860_ = _02859_ | _02858_;
  assign _02861_ = sel_oi_one_hot_i[126] & i[233];
  assign _02862_ = sel_oi_one_hot_i[127] & i[249];
  assign _02863_ = _02862_ | _02861_;
  assign _02864_ = _02863_ | _02860_;
  assign _02865_ = _02864_ | _02857_;
  assign o[121] = _02865_ | _02850_;
  assign _02866_ = sel_oi_one_hot_i[112] & i[8];
  assign _02867_ = sel_oi_one_hot_i[113] & i[24];
  assign _02868_ = _02867_ | _02866_;
  assign _02869_ = sel_oi_one_hot_i[114] & i[40];
  assign _02870_ = sel_oi_one_hot_i[115] & i[56];
  assign _02871_ = _02870_ | _02869_;
  assign _02872_ = _02871_ | _02868_;
  assign _02873_ = sel_oi_one_hot_i[116] & i[72];
  assign _02874_ = sel_oi_one_hot_i[117] & i[88];
  assign _02875_ = _02874_ | _02873_;
  assign _02876_ = sel_oi_one_hot_i[118] & i[104];
  assign _02877_ = sel_oi_one_hot_i[119] & i[120];
  assign _02878_ = _02877_ | _02876_;
  assign _02879_ = _02878_ | _02875_;
  assign _02880_ = _02879_ | _02872_;
  assign _02881_ = sel_oi_one_hot_i[120] & i[136];
  assign _02882_ = sel_oi_one_hot_i[121] & i[152];
  assign _02883_ = _02882_ | _02881_;
  assign _02884_ = sel_oi_one_hot_i[122] & i[168];
  assign _02885_ = sel_oi_one_hot_i[123] & i[184];
  assign _02886_ = _02885_ | _02884_;
  assign _02887_ = _02886_ | _02883_;
  assign _02888_ = sel_oi_one_hot_i[124] & i[200];
  assign _02889_ = sel_oi_one_hot_i[125] & i[216];
  assign _02890_ = _02889_ | _02888_;
  assign _02891_ = sel_oi_one_hot_i[126] & i[232];
  assign _02892_ = sel_oi_one_hot_i[127] & i[248];
  assign _02893_ = _02892_ | _02891_;
  assign _02894_ = _02893_ | _02890_;
  assign _02895_ = _02894_ | _02887_;
  assign o[120] = _02895_ | _02880_;
  assign _02896_ = sel_oi_one_hot_i[112] & i[7];
  assign _02897_ = sel_oi_one_hot_i[113] & i[23];
  assign _02898_ = _02897_ | _02896_;
  assign _02899_ = sel_oi_one_hot_i[114] & i[39];
  assign _02900_ = sel_oi_one_hot_i[115] & i[55];
  assign _02901_ = _02900_ | _02899_;
  assign _02902_ = _02901_ | _02898_;
  assign _02903_ = sel_oi_one_hot_i[116] & i[71];
  assign _02904_ = sel_oi_one_hot_i[117] & i[87];
  assign _02905_ = _02904_ | _02903_;
  assign _02906_ = sel_oi_one_hot_i[118] & i[103];
  assign _02907_ = sel_oi_one_hot_i[119] & i[119];
  assign _02908_ = _02907_ | _02906_;
  assign _02909_ = _02908_ | _02905_;
  assign _02910_ = _02909_ | _02902_;
  assign _02911_ = sel_oi_one_hot_i[120] & i[135];
  assign _02912_ = sel_oi_one_hot_i[121] & i[151];
  assign _02913_ = _02912_ | _02911_;
  assign _02914_ = sel_oi_one_hot_i[122] & i[167];
  assign _02915_ = sel_oi_one_hot_i[123] & i[183];
  assign _02916_ = _02915_ | _02914_;
  assign _02917_ = _02916_ | _02913_;
  assign _02918_ = sel_oi_one_hot_i[124] & i[199];
  assign _02919_ = sel_oi_one_hot_i[125] & i[215];
  assign _02920_ = _02919_ | _02918_;
  assign _02921_ = sel_oi_one_hot_i[126] & i[231];
  assign _02922_ = sel_oi_one_hot_i[127] & i[247];
  assign _02923_ = _02922_ | _02921_;
  assign _02924_ = _02923_ | _02920_;
  assign _02925_ = _02924_ | _02917_;
  assign o[119] = _02925_ | _02910_;
  assign _02926_ = sel_oi_one_hot_i[112] & i[6];
  assign _02927_ = sel_oi_one_hot_i[113] & i[22];
  assign _02928_ = _02927_ | _02926_;
  assign _02929_ = sel_oi_one_hot_i[114] & i[38];
  assign _02930_ = sel_oi_one_hot_i[115] & i[54];
  assign _02931_ = _02930_ | _02929_;
  assign _02932_ = _02931_ | _02928_;
  assign _02933_ = sel_oi_one_hot_i[116] & i[70];
  assign _02934_ = sel_oi_one_hot_i[117] & i[86];
  assign _02935_ = _02934_ | _02933_;
  assign _02936_ = sel_oi_one_hot_i[118] & i[102];
  assign _02937_ = sel_oi_one_hot_i[119] & i[118];
  assign _02938_ = _02937_ | _02936_;
  assign _02939_ = _02938_ | _02935_;
  assign _02940_ = _02939_ | _02932_;
  assign _02941_ = sel_oi_one_hot_i[120] & i[134];
  assign _02942_ = sel_oi_one_hot_i[121] & i[150];
  assign _02943_ = _02942_ | _02941_;
  assign _02944_ = sel_oi_one_hot_i[122] & i[166];
  assign _02945_ = sel_oi_one_hot_i[123] & i[182];
  assign _02946_ = _02945_ | _02944_;
  assign _02947_ = _02946_ | _02943_;
  assign _02948_ = sel_oi_one_hot_i[124] & i[198];
  assign _02949_ = sel_oi_one_hot_i[125] & i[214];
  assign _02950_ = _02949_ | _02948_;
  assign _02951_ = sel_oi_one_hot_i[126] & i[230];
  assign _02952_ = sel_oi_one_hot_i[127] & i[246];
  assign _02953_ = _02952_ | _02951_;
  assign _02954_ = _02953_ | _02950_;
  assign _02955_ = _02954_ | _02947_;
  assign o[118] = _02955_ | _02940_;
  assign _02956_ = sel_oi_one_hot_i[112] & i[5];
  assign _02957_ = sel_oi_one_hot_i[113] & i[21];
  assign _02958_ = _02957_ | _02956_;
  assign _02959_ = sel_oi_one_hot_i[114] & i[37];
  assign _02960_ = sel_oi_one_hot_i[115] & i[53];
  assign _02961_ = _02960_ | _02959_;
  assign _02962_ = _02961_ | _02958_;
  assign _02963_ = sel_oi_one_hot_i[116] & i[69];
  assign _02964_ = sel_oi_one_hot_i[117] & i[85];
  assign _02965_ = _02964_ | _02963_;
  assign _02966_ = sel_oi_one_hot_i[118] & i[101];
  assign _02967_ = sel_oi_one_hot_i[119] & i[117];
  assign _02968_ = _02967_ | _02966_;
  assign _02969_ = _02968_ | _02965_;
  assign _02970_ = _02969_ | _02962_;
  assign _02971_ = sel_oi_one_hot_i[120] & i[133];
  assign _02972_ = sel_oi_one_hot_i[121] & i[149];
  assign _02973_ = _02972_ | _02971_;
  assign _02974_ = sel_oi_one_hot_i[122] & i[165];
  assign _02975_ = sel_oi_one_hot_i[123] & i[181];
  assign _02976_ = _02975_ | _02974_;
  assign _02977_ = _02976_ | _02973_;
  assign _02978_ = sel_oi_one_hot_i[124] & i[197];
  assign _02979_ = sel_oi_one_hot_i[125] & i[213];
  assign _02980_ = _02979_ | _02978_;
  assign _02981_ = sel_oi_one_hot_i[126] & i[229];
  assign _02982_ = sel_oi_one_hot_i[127] & i[245];
  assign _02983_ = _02982_ | _02981_;
  assign _02984_ = _02983_ | _02980_;
  assign _02985_ = _02984_ | _02977_;
  assign o[117] = _02985_ | _02970_;
  assign _02986_ = sel_oi_one_hot_i[112] & i[4];
  assign _02987_ = sel_oi_one_hot_i[113] & i[20];
  assign _02988_ = _02987_ | _02986_;
  assign _02989_ = sel_oi_one_hot_i[114] & i[36];
  assign _02990_ = sel_oi_one_hot_i[115] & i[52];
  assign _02991_ = _02990_ | _02989_;
  assign _02992_ = _02991_ | _02988_;
  assign _02993_ = sel_oi_one_hot_i[116] & i[68];
  assign _02994_ = sel_oi_one_hot_i[117] & i[84];
  assign _02995_ = _02994_ | _02993_;
  assign _02996_ = sel_oi_one_hot_i[118] & i[100];
  assign _02997_ = sel_oi_one_hot_i[119] & i[116];
  assign _02998_ = _02997_ | _02996_;
  assign _02999_ = _02998_ | _02995_;
  assign _03000_ = _02999_ | _02992_;
  assign _03001_ = sel_oi_one_hot_i[120] & i[132];
  assign _03002_ = sel_oi_one_hot_i[121] & i[148];
  assign _03003_ = _03002_ | _03001_;
  assign _03004_ = sel_oi_one_hot_i[122] & i[164];
  assign _03005_ = sel_oi_one_hot_i[123] & i[180];
  assign _03006_ = _03005_ | _03004_;
  assign _03007_ = _03006_ | _03003_;
  assign _03008_ = sel_oi_one_hot_i[124] & i[196];
  assign _03009_ = sel_oi_one_hot_i[125] & i[212];
  assign _03010_ = _03009_ | _03008_;
  assign _03011_ = sel_oi_one_hot_i[126] & i[228];
  assign _03012_ = sel_oi_one_hot_i[127] & i[244];
  assign _03013_ = _03012_ | _03011_;
  assign _03014_ = _03013_ | _03010_;
  assign _03015_ = _03014_ | _03007_;
  assign o[116] = _03015_ | _03000_;
  assign _03016_ = sel_oi_one_hot_i[112] & i[3];
  assign _03017_ = sel_oi_one_hot_i[113] & i[19];
  assign _03018_ = _03017_ | _03016_;
  assign _03019_ = sel_oi_one_hot_i[114] & i[35];
  assign _03020_ = sel_oi_one_hot_i[115] & i[51];
  assign _03021_ = _03020_ | _03019_;
  assign _03022_ = _03021_ | _03018_;
  assign _03023_ = sel_oi_one_hot_i[116] & i[67];
  assign _03024_ = sel_oi_one_hot_i[117] & i[83];
  assign _03025_ = _03024_ | _03023_;
  assign _03026_ = sel_oi_one_hot_i[118] & i[99];
  assign _03027_ = sel_oi_one_hot_i[119] & i[115];
  assign _03028_ = _03027_ | _03026_;
  assign _03029_ = _03028_ | _03025_;
  assign _03030_ = _03029_ | _03022_;
  assign _03031_ = sel_oi_one_hot_i[120] & i[131];
  assign _03032_ = sel_oi_one_hot_i[121] & i[147];
  assign _03033_ = _03032_ | _03031_;
  assign _03034_ = sel_oi_one_hot_i[122] & i[163];
  assign _03035_ = sel_oi_one_hot_i[123] & i[179];
  assign _03036_ = _03035_ | _03034_;
  assign _03037_ = _03036_ | _03033_;
  assign _03038_ = sel_oi_one_hot_i[124] & i[195];
  assign _03039_ = sel_oi_one_hot_i[125] & i[211];
  assign _03040_ = _03039_ | _03038_;
  assign _03041_ = sel_oi_one_hot_i[126] & i[227];
  assign _03042_ = sel_oi_one_hot_i[127] & i[243];
  assign _03043_ = _03042_ | _03041_;
  assign _03044_ = _03043_ | _03040_;
  assign _03045_ = _03044_ | _03037_;
  assign o[115] = _03045_ | _03030_;
  assign _03046_ = sel_oi_one_hot_i[112] & i[2];
  assign _03047_ = sel_oi_one_hot_i[113] & i[18];
  assign _03048_ = _03047_ | _03046_;
  assign _03049_ = sel_oi_one_hot_i[114] & i[34];
  assign _03050_ = sel_oi_one_hot_i[115] & i[50];
  assign _03051_ = _03050_ | _03049_;
  assign _03052_ = _03051_ | _03048_;
  assign _03053_ = sel_oi_one_hot_i[116] & i[66];
  assign _03054_ = sel_oi_one_hot_i[117] & i[82];
  assign _03055_ = _03054_ | _03053_;
  assign _03056_ = sel_oi_one_hot_i[118] & i[98];
  assign _03057_ = sel_oi_one_hot_i[119] & i[114];
  assign _03058_ = _03057_ | _03056_;
  assign _03059_ = _03058_ | _03055_;
  assign _03060_ = _03059_ | _03052_;
  assign _03061_ = sel_oi_one_hot_i[120] & i[130];
  assign _03062_ = sel_oi_one_hot_i[121] & i[146];
  assign _03063_ = _03062_ | _03061_;
  assign _03064_ = sel_oi_one_hot_i[122] & i[162];
  assign _03065_ = sel_oi_one_hot_i[123] & i[178];
  assign _03066_ = _03065_ | _03064_;
  assign _03067_ = _03066_ | _03063_;
  assign _03068_ = sel_oi_one_hot_i[124] & i[194];
  assign _03069_ = sel_oi_one_hot_i[125] & i[210];
  assign _03070_ = _03069_ | _03068_;
  assign _03071_ = sel_oi_one_hot_i[126] & i[226];
  assign _03072_ = sel_oi_one_hot_i[127] & i[242];
  assign _03073_ = _03072_ | _03071_;
  assign _03074_ = _03073_ | _03070_;
  assign _03075_ = _03074_ | _03067_;
  assign o[114] = _03075_ | _03060_;
  assign _03076_ = sel_oi_one_hot_i[112] & i[1];
  assign _03077_ = sel_oi_one_hot_i[113] & i[17];
  assign _03078_ = _03077_ | _03076_;
  assign _03079_ = sel_oi_one_hot_i[114] & i[33];
  assign _03080_ = sel_oi_one_hot_i[115] & i[49];
  assign _03081_ = _03080_ | _03079_;
  assign _03082_ = _03081_ | _03078_;
  assign _03083_ = sel_oi_one_hot_i[116] & i[65];
  assign _03084_ = sel_oi_one_hot_i[117] & i[81];
  assign _03085_ = _03084_ | _03083_;
  assign _03086_ = sel_oi_one_hot_i[118] & i[97];
  assign _03087_ = sel_oi_one_hot_i[119] & i[113];
  assign _03088_ = _03087_ | _03086_;
  assign _03089_ = _03088_ | _03085_;
  assign _03090_ = _03089_ | _03082_;
  assign _03091_ = sel_oi_one_hot_i[120] & i[129];
  assign _03092_ = sel_oi_one_hot_i[121] & i[145];
  assign _03093_ = _03092_ | _03091_;
  assign _03094_ = sel_oi_one_hot_i[122] & i[161];
  assign _03095_ = sel_oi_one_hot_i[123] & i[177];
  assign _03096_ = _03095_ | _03094_;
  assign _03097_ = _03096_ | _03093_;
  assign _03098_ = sel_oi_one_hot_i[124] & i[193];
  assign _03099_ = sel_oi_one_hot_i[125] & i[209];
  assign _03100_ = _03099_ | _03098_;
  assign _03101_ = sel_oi_one_hot_i[126] & i[225];
  assign _03102_ = sel_oi_one_hot_i[127] & i[241];
  assign _03103_ = _03102_ | _03101_;
  assign _03104_ = _03103_ | _03100_;
  assign _03105_ = _03104_ | _03097_;
  assign o[113] = _03105_ | _03090_;
  assign _03106_ = sel_oi_one_hot_i[112] & i[0];
  assign _03107_ = sel_oi_one_hot_i[113] & i[16];
  assign _03108_ = _03107_ | _03106_;
  assign _03109_ = sel_oi_one_hot_i[114] & i[32];
  assign _03110_ = sel_oi_one_hot_i[115] & i[48];
  assign _03111_ = _03110_ | _03109_;
  assign _03112_ = _03111_ | _03108_;
  assign _03113_ = sel_oi_one_hot_i[116] & i[64];
  assign _03114_ = sel_oi_one_hot_i[117] & i[80];
  assign _03115_ = _03114_ | _03113_;
  assign _03116_ = sel_oi_one_hot_i[118] & i[96];
  assign _03117_ = sel_oi_one_hot_i[119] & i[112];
  assign _03118_ = _03117_ | _03116_;
  assign _03119_ = _03118_ | _03115_;
  assign _03120_ = _03119_ | _03112_;
  assign _03121_ = sel_oi_one_hot_i[120] & i[128];
  assign _03122_ = sel_oi_one_hot_i[121] & i[144];
  assign _03123_ = _03122_ | _03121_;
  assign _03124_ = sel_oi_one_hot_i[122] & i[160];
  assign _03125_ = sel_oi_one_hot_i[123] & i[176];
  assign _03126_ = _03125_ | _03124_;
  assign _03127_ = _03126_ | _03123_;
  assign _03128_ = sel_oi_one_hot_i[124] & i[192];
  assign _03129_ = sel_oi_one_hot_i[125] & i[208];
  assign _03130_ = _03129_ | _03128_;
  assign _03131_ = sel_oi_one_hot_i[126] & i[224];
  assign _03132_ = sel_oi_one_hot_i[127] & i[240];
  assign _03133_ = _03132_ | _03131_;
  assign _03134_ = _03133_ | _03130_;
  assign _03135_ = _03134_ | _03127_;
  assign o[112] = _03135_ | _03120_;
  assign _03136_ = sel_oi_one_hot_i[128] & i[15];
  assign _03137_ = sel_oi_one_hot_i[129] & i[31];
  assign _03138_ = _03137_ | _03136_;
  assign _03139_ = sel_oi_one_hot_i[130] & i[47];
  assign _03140_ = sel_oi_one_hot_i[131] & i[63];
  assign _03141_ = _03140_ | _03139_;
  assign _03142_ = _03141_ | _03138_;
  assign _03143_ = sel_oi_one_hot_i[132] & i[79];
  assign _03144_ = sel_oi_one_hot_i[133] & i[95];
  assign _03145_ = _03144_ | _03143_;
  assign _03146_ = sel_oi_one_hot_i[134] & i[111];
  assign _03147_ = sel_oi_one_hot_i[135] & i[127];
  assign _03148_ = _03147_ | _03146_;
  assign _03149_ = _03148_ | _03145_;
  assign _03150_ = _03149_ | _03142_;
  assign _03151_ = sel_oi_one_hot_i[136] & i[143];
  assign _03152_ = sel_oi_one_hot_i[137] & i[159];
  assign _03153_ = _03152_ | _03151_;
  assign _03154_ = sel_oi_one_hot_i[138] & i[175];
  assign _03155_ = sel_oi_one_hot_i[139] & i[191];
  assign _03156_ = _03155_ | _03154_;
  assign _03157_ = _03156_ | _03153_;
  assign _03158_ = sel_oi_one_hot_i[140] & i[207];
  assign _03159_ = sel_oi_one_hot_i[141] & i[223];
  assign _03160_ = _03159_ | _03158_;
  assign _03161_ = sel_oi_one_hot_i[142] & i[239];
  assign _03162_ = sel_oi_one_hot_i[143] & i[255];
  assign _03163_ = _03162_ | _03161_;
  assign _03164_ = _03163_ | _03160_;
  assign _03165_ = _03164_ | _03157_;
  assign o[143] = _03165_ | _03150_;
  assign _03166_ = sel_oi_one_hot_i[128] & i[14];
  assign _03167_ = sel_oi_one_hot_i[129] & i[30];
  assign _03168_ = _03167_ | _03166_;
  assign _03169_ = sel_oi_one_hot_i[130] & i[46];
  assign _03170_ = sel_oi_one_hot_i[131] & i[62];
  assign _03171_ = _03170_ | _03169_;
  assign _03172_ = _03171_ | _03168_;
  assign _03173_ = sel_oi_one_hot_i[132] & i[78];
  assign _03174_ = sel_oi_one_hot_i[133] & i[94];
  assign _03175_ = _03174_ | _03173_;
  assign _03176_ = sel_oi_one_hot_i[134] & i[110];
  assign _03177_ = sel_oi_one_hot_i[135] & i[126];
  assign _03178_ = _03177_ | _03176_;
  assign _03179_ = _03178_ | _03175_;
  assign _03180_ = _03179_ | _03172_;
  assign _03181_ = sel_oi_one_hot_i[136] & i[142];
  assign _03182_ = sel_oi_one_hot_i[137] & i[158];
  assign _03183_ = _03182_ | _03181_;
  assign _03184_ = sel_oi_one_hot_i[138] & i[174];
  assign _03185_ = sel_oi_one_hot_i[139] & i[190];
  assign _03186_ = _03185_ | _03184_;
  assign _03187_ = _03186_ | _03183_;
  assign _03188_ = sel_oi_one_hot_i[140] & i[206];
  assign _03189_ = sel_oi_one_hot_i[141] & i[222];
  assign _03190_ = _03189_ | _03188_;
  assign _03191_ = sel_oi_one_hot_i[142] & i[238];
  assign _03192_ = sel_oi_one_hot_i[143] & i[254];
  assign _03193_ = _03192_ | _03191_;
  assign _03194_ = _03193_ | _03190_;
  assign _03195_ = _03194_ | _03187_;
  assign o[142] = _03195_ | _03180_;
  assign _03196_ = sel_oi_one_hot_i[128] & i[13];
  assign _03197_ = sel_oi_one_hot_i[129] & i[29];
  assign _03198_ = _03197_ | _03196_;
  assign _03199_ = sel_oi_one_hot_i[130] & i[45];
  assign _03200_ = sel_oi_one_hot_i[131] & i[61];
  assign _03201_ = _03200_ | _03199_;
  assign _03202_ = _03201_ | _03198_;
  assign _03203_ = sel_oi_one_hot_i[132] & i[77];
  assign _03204_ = sel_oi_one_hot_i[133] & i[93];
  assign _03205_ = _03204_ | _03203_;
  assign _03206_ = sel_oi_one_hot_i[134] & i[109];
  assign _03207_ = sel_oi_one_hot_i[135] & i[125];
  assign _03208_ = _03207_ | _03206_;
  assign _03209_ = _03208_ | _03205_;
  assign _03210_ = _03209_ | _03202_;
  assign _03211_ = sel_oi_one_hot_i[136] & i[141];
  assign _03212_ = sel_oi_one_hot_i[137] & i[157];
  assign _03213_ = _03212_ | _03211_;
  assign _03214_ = sel_oi_one_hot_i[138] & i[173];
  assign _03215_ = sel_oi_one_hot_i[139] & i[189];
  assign _03216_ = _03215_ | _03214_;
  assign _03217_ = _03216_ | _03213_;
  assign _03218_ = sel_oi_one_hot_i[140] & i[205];
  assign _03219_ = sel_oi_one_hot_i[141] & i[221];
  assign _03220_ = _03219_ | _03218_;
  assign _03221_ = sel_oi_one_hot_i[142] & i[237];
  assign _03222_ = sel_oi_one_hot_i[143] & i[253];
  assign _03223_ = _03222_ | _03221_;
  assign _03224_ = _03223_ | _03220_;
  assign _03225_ = _03224_ | _03217_;
  assign o[141] = _03225_ | _03210_;
  assign _03226_ = sel_oi_one_hot_i[128] & i[12];
  assign _03227_ = sel_oi_one_hot_i[129] & i[28];
  assign _03228_ = _03227_ | _03226_;
  assign _03229_ = sel_oi_one_hot_i[130] & i[44];
  assign _03230_ = sel_oi_one_hot_i[131] & i[60];
  assign _03231_ = _03230_ | _03229_;
  assign _03232_ = _03231_ | _03228_;
  assign _03233_ = sel_oi_one_hot_i[132] & i[76];
  assign _03234_ = sel_oi_one_hot_i[133] & i[92];
  assign _03235_ = _03234_ | _03233_;
  assign _03236_ = sel_oi_one_hot_i[134] & i[108];
  assign _03237_ = sel_oi_one_hot_i[135] & i[124];
  assign _03238_ = _03237_ | _03236_;
  assign _03239_ = _03238_ | _03235_;
  assign _03240_ = _03239_ | _03232_;
  assign _03241_ = sel_oi_one_hot_i[136] & i[140];
  assign _03242_ = sel_oi_one_hot_i[137] & i[156];
  assign _03243_ = _03242_ | _03241_;
  assign _03244_ = sel_oi_one_hot_i[138] & i[172];
  assign _03245_ = sel_oi_one_hot_i[139] & i[188];
  assign _03246_ = _03245_ | _03244_;
  assign _03247_ = _03246_ | _03243_;
  assign _03248_ = sel_oi_one_hot_i[140] & i[204];
  assign _03249_ = sel_oi_one_hot_i[141] & i[220];
  assign _03250_ = _03249_ | _03248_;
  assign _03251_ = sel_oi_one_hot_i[142] & i[236];
  assign _03252_ = sel_oi_one_hot_i[143] & i[252];
  assign _03253_ = _03252_ | _03251_;
  assign _03254_ = _03253_ | _03250_;
  assign _03255_ = _03254_ | _03247_;
  assign o[140] = _03255_ | _03240_;
  assign _03256_ = sel_oi_one_hot_i[128] & i[11];
  assign _03257_ = sel_oi_one_hot_i[129] & i[27];
  assign _03258_ = _03257_ | _03256_;
  assign _03259_ = sel_oi_one_hot_i[130] & i[43];
  assign _03260_ = sel_oi_one_hot_i[131] & i[59];
  assign _03261_ = _03260_ | _03259_;
  assign _03262_ = _03261_ | _03258_;
  assign _03263_ = sel_oi_one_hot_i[132] & i[75];
  assign _03264_ = sel_oi_one_hot_i[133] & i[91];
  assign _03265_ = _03264_ | _03263_;
  assign _03266_ = sel_oi_one_hot_i[134] & i[107];
  assign _03267_ = sel_oi_one_hot_i[135] & i[123];
  assign _03268_ = _03267_ | _03266_;
  assign _03269_ = _03268_ | _03265_;
  assign _03270_ = _03269_ | _03262_;
  assign _03271_ = sel_oi_one_hot_i[136] & i[139];
  assign _03272_ = sel_oi_one_hot_i[137] & i[155];
  assign _03273_ = _03272_ | _03271_;
  assign _03274_ = sel_oi_one_hot_i[138] & i[171];
  assign _03275_ = sel_oi_one_hot_i[139] & i[187];
  assign _03276_ = _03275_ | _03274_;
  assign _03277_ = _03276_ | _03273_;
  assign _03278_ = sel_oi_one_hot_i[140] & i[203];
  assign _03279_ = sel_oi_one_hot_i[141] & i[219];
  assign _03280_ = _03279_ | _03278_;
  assign _03281_ = sel_oi_one_hot_i[142] & i[235];
  assign _03282_ = sel_oi_one_hot_i[143] & i[251];
  assign _03283_ = _03282_ | _03281_;
  assign _03284_ = _03283_ | _03280_;
  assign _03285_ = _03284_ | _03277_;
  assign o[139] = _03285_ | _03270_;
  assign _03286_ = sel_oi_one_hot_i[128] & i[10];
  assign _03287_ = sel_oi_one_hot_i[129] & i[26];
  assign _03288_ = _03287_ | _03286_;
  assign _03289_ = sel_oi_one_hot_i[130] & i[42];
  assign _03290_ = sel_oi_one_hot_i[131] & i[58];
  assign _03291_ = _03290_ | _03289_;
  assign _03292_ = _03291_ | _03288_;
  assign _03293_ = sel_oi_one_hot_i[132] & i[74];
  assign _03294_ = sel_oi_one_hot_i[133] & i[90];
  assign _03295_ = _03294_ | _03293_;
  assign _03296_ = sel_oi_one_hot_i[134] & i[106];
  assign _03297_ = sel_oi_one_hot_i[135] & i[122];
  assign _03298_ = _03297_ | _03296_;
  assign _03299_ = _03298_ | _03295_;
  assign _03300_ = _03299_ | _03292_;
  assign _03301_ = sel_oi_one_hot_i[136] & i[138];
  assign _03302_ = sel_oi_one_hot_i[137] & i[154];
  assign _03303_ = _03302_ | _03301_;
  assign _03304_ = sel_oi_one_hot_i[138] & i[170];
  assign _03305_ = sel_oi_one_hot_i[139] & i[186];
  assign _03306_ = _03305_ | _03304_;
  assign _03307_ = _03306_ | _03303_;
  assign _03308_ = sel_oi_one_hot_i[140] & i[202];
  assign _03309_ = sel_oi_one_hot_i[141] & i[218];
  assign _03310_ = _03309_ | _03308_;
  assign _03311_ = sel_oi_one_hot_i[142] & i[234];
  assign _03312_ = sel_oi_one_hot_i[143] & i[250];
  assign _03313_ = _03312_ | _03311_;
  assign _03314_ = _03313_ | _03310_;
  assign _03315_ = _03314_ | _03307_;
  assign o[138] = _03315_ | _03300_;
  assign _03316_ = sel_oi_one_hot_i[128] & i[9];
  assign _03317_ = sel_oi_one_hot_i[129] & i[25];
  assign _03318_ = _03317_ | _03316_;
  assign _03319_ = sel_oi_one_hot_i[130] & i[41];
  assign _03320_ = sel_oi_one_hot_i[131] & i[57];
  assign _03321_ = _03320_ | _03319_;
  assign _03322_ = _03321_ | _03318_;
  assign _03323_ = sel_oi_one_hot_i[132] & i[73];
  assign _03324_ = sel_oi_one_hot_i[133] & i[89];
  assign _03325_ = _03324_ | _03323_;
  assign _03326_ = sel_oi_one_hot_i[134] & i[105];
  assign _03327_ = sel_oi_one_hot_i[135] & i[121];
  assign _03328_ = _03327_ | _03326_;
  assign _03329_ = _03328_ | _03325_;
  assign _03330_ = _03329_ | _03322_;
  assign _03331_ = sel_oi_one_hot_i[136] & i[137];
  assign _03332_ = sel_oi_one_hot_i[137] & i[153];
  assign _03333_ = _03332_ | _03331_;
  assign _03334_ = sel_oi_one_hot_i[138] & i[169];
  assign _03335_ = sel_oi_one_hot_i[139] & i[185];
  assign _03336_ = _03335_ | _03334_;
  assign _03337_ = _03336_ | _03333_;
  assign _03338_ = sel_oi_one_hot_i[140] & i[201];
  assign _03339_ = sel_oi_one_hot_i[141] & i[217];
  assign _03340_ = _03339_ | _03338_;
  assign _03341_ = sel_oi_one_hot_i[142] & i[233];
  assign _03342_ = sel_oi_one_hot_i[143] & i[249];
  assign _03343_ = _03342_ | _03341_;
  assign _03344_ = _03343_ | _03340_;
  assign _03345_ = _03344_ | _03337_;
  assign o[137] = _03345_ | _03330_;
  assign _03346_ = sel_oi_one_hot_i[128] & i[8];
  assign _03347_ = sel_oi_one_hot_i[129] & i[24];
  assign _03348_ = _03347_ | _03346_;
  assign _03349_ = sel_oi_one_hot_i[130] & i[40];
  assign _03350_ = sel_oi_one_hot_i[131] & i[56];
  assign _03351_ = _03350_ | _03349_;
  assign _03352_ = _03351_ | _03348_;
  assign _03353_ = sel_oi_one_hot_i[132] & i[72];
  assign _03354_ = sel_oi_one_hot_i[133] & i[88];
  assign _03355_ = _03354_ | _03353_;
  assign _03356_ = sel_oi_one_hot_i[134] & i[104];
  assign _03357_ = sel_oi_one_hot_i[135] & i[120];
  assign _03358_ = _03357_ | _03356_;
  assign _03359_ = _03358_ | _03355_;
  assign _03360_ = _03359_ | _03352_;
  assign _03361_ = sel_oi_one_hot_i[136] & i[136];
  assign _03362_ = sel_oi_one_hot_i[137] & i[152];
  assign _03363_ = _03362_ | _03361_;
  assign _03364_ = sel_oi_one_hot_i[138] & i[168];
  assign _03365_ = sel_oi_one_hot_i[139] & i[184];
  assign _03366_ = _03365_ | _03364_;
  assign _03367_ = _03366_ | _03363_;
  assign _03368_ = sel_oi_one_hot_i[140] & i[200];
  assign _03369_ = sel_oi_one_hot_i[141] & i[216];
  assign _03370_ = _03369_ | _03368_;
  assign _03371_ = sel_oi_one_hot_i[142] & i[232];
  assign _03372_ = sel_oi_one_hot_i[143] & i[248];
  assign _03373_ = _03372_ | _03371_;
  assign _03374_ = _03373_ | _03370_;
  assign _03375_ = _03374_ | _03367_;
  assign o[136] = _03375_ | _03360_;
  assign _03376_ = sel_oi_one_hot_i[128] & i[7];
  assign _03377_ = sel_oi_one_hot_i[129] & i[23];
  assign _03378_ = _03377_ | _03376_;
  assign _03379_ = sel_oi_one_hot_i[130] & i[39];
  assign _03380_ = sel_oi_one_hot_i[131] & i[55];
  assign _03381_ = _03380_ | _03379_;
  assign _03382_ = _03381_ | _03378_;
  assign _03383_ = sel_oi_one_hot_i[132] & i[71];
  assign _03384_ = sel_oi_one_hot_i[133] & i[87];
  assign _03385_ = _03384_ | _03383_;
  assign _03386_ = sel_oi_one_hot_i[134] & i[103];
  assign _03387_ = sel_oi_one_hot_i[135] & i[119];
  assign _03388_ = _03387_ | _03386_;
  assign _03389_ = _03388_ | _03385_;
  assign _03390_ = _03389_ | _03382_;
  assign _03391_ = sel_oi_one_hot_i[136] & i[135];
  assign _03392_ = sel_oi_one_hot_i[137] & i[151];
  assign _03393_ = _03392_ | _03391_;
  assign _03394_ = sel_oi_one_hot_i[138] & i[167];
  assign _03395_ = sel_oi_one_hot_i[139] & i[183];
  assign _03396_ = _03395_ | _03394_;
  assign _03397_ = _03396_ | _03393_;
  assign _03398_ = sel_oi_one_hot_i[140] & i[199];
  assign _03399_ = sel_oi_one_hot_i[141] & i[215];
  assign _03400_ = _03399_ | _03398_;
  assign _03401_ = sel_oi_one_hot_i[142] & i[231];
  assign _03402_ = sel_oi_one_hot_i[143] & i[247];
  assign _03403_ = _03402_ | _03401_;
  assign _03404_ = _03403_ | _03400_;
  assign _03405_ = _03404_ | _03397_;
  assign o[135] = _03405_ | _03390_;
  assign _03406_ = sel_oi_one_hot_i[128] & i[6];
  assign _03407_ = sel_oi_one_hot_i[129] & i[22];
  assign _03408_ = _03407_ | _03406_;
  assign _03409_ = sel_oi_one_hot_i[130] & i[38];
  assign _03410_ = sel_oi_one_hot_i[131] & i[54];
  assign _03411_ = _03410_ | _03409_;
  assign _03412_ = _03411_ | _03408_;
  assign _03413_ = sel_oi_one_hot_i[132] & i[70];
  assign _03414_ = sel_oi_one_hot_i[133] & i[86];
  assign _03415_ = _03414_ | _03413_;
  assign _03416_ = sel_oi_one_hot_i[134] & i[102];
  assign _03417_ = sel_oi_one_hot_i[135] & i[118];
  assign _03418_ = _03417_ | _03416_;
  assign _03419_ = _03418_ | _03415_;
  assign _03420_ = _03419_ | _03412_;
  assign _03421_ = sel_oi_one_hot_i[136] & i[134];
  assign _03422_ = sel_oi_one_hot_i[137] & i[150];
  assign _03423_ = _03422_ | _03421_;
  assign _03424_ = sel_oi_one_hot_i[138] & i[166];
  assign _03425_ = sel_oi_one_hot_i[139] & i[182];
  assign _03426_ = _03425_ | _03424_;
  assign _03427_ = _03426_ | _03423_;
  assign _03428_ = sel_oi_one_hot_i[140] & i[198];
  assign _03429_ = sel_oi_one_hot_i[141] & i[214];
  assign _03430_ = _03429_ | _03428_;
  assign _03431_ = sel_oi_one_hot_i[142] & i[230];
  assign _03432_ = sel_oi_one_hot_i[143] & i[246];
  assign _03433_ = _03432_ | _03431_;
  assign _03434_ = _03433_ | _03430_;
  assign _03435_ = _03434_ | _03427_;
  assign o[134] = _03435_ | _03420_;
  assign _03436_ = sel_oi_one_hot_i[128] & i[5];
  assign _03437_ = sel_oi_one_hot_i[129] & i[21];
  assign _03438_ = _03437_ | _03436_;
  assign _03439_ = sel_oi_one_hot_i[130] & i[37];
  assign _03440_ = sel_oi_one_hot_i[131] & i[53];
  assign _03441_ = _03440_ | _03439_;
  assign _03442_ = _03441_ | _03438_;
  assign _03443_ = sel_oi_one_hot_i[132] & i[69];
  assign _03444_ = sel_oi_one_hot_i[133] & i[85];
  assign _03445_ = _03444_ | _03443_;
  assign _03446_ = sel_oi_one_hot_i[134] & i[101];
  assign _03447_ = sel_oi_one_hot_i[135] & i[117];
  assign _03448_ = _03447_ | _03446_;
  assign _03449_ = _03448_ | _03445_;
  assign _03450_ = _03449_ | _03442_;
  assign _03451_ = sel_oi_one_hot_i[136] & i[133];
  assign _03452_ = sel_oi_one_hot_i[137] & i[149];
  assign _03453_ = _03452_ | _03451_;
  assign _03454_ = sel_oi_one_hot_i[138] & i[165];
  assign _03455_ = sel_oi_one_hot_i[139] & i[181];
  assign _03456_ = _03455_ | _03454_;
  assign _03457_ = _03456_ | _03453_;
  assign _03458_ = sel_oi_one_hot_i[140] & i[197];
  assign _03459_ = sel_oi_one_hot_i[141] & i[213];
  assign _03460_ = _03459_ | _03458_;
  assign _03461_ = sel_oi_one_hot_i[142] & i[229];
  assign _03462_ = sel_oi_one_hot_i[143] & i[245];
  assign _03463_ = _03462_ | _03461_;
  assign _03464_ = _03463_ | _03460_;
  assign _03465_ = _03464_ | _03457_;
  assign o[133] = _03465_ | _03450_;
  assign _03466_ = sel_oi_one_hot_i[128] & i[4];
  assign _03467_ = sel_oi_one_hot_i[129] & i[20];
  assign _03468_ = _03467_ | _03466_;
  assign _03469_ = sel_oi_one_hot_i[130] & i[36];
  assign _03470_ = sel_oi_one_hot_i[131] & i[52];
  assign _03471_ = _03470_ | _03469_;
  assign _03472_ = _03471_ | _03468_;
  assign _03473_ = sel_oi_one_hot_i[132] & i[68];
  assign _03474_ = sel_oi_one_hot_i[133] & i[84];
  assign _03475_ = _03474_ | _03473_;
  assign _03476_ = sel_oi_one_hot_i[134] & i[100];
  assign _03477_ = sel_oi_one_hot_i[135] & i[116];
  assign _03478_ = _03477_ | _03476_;
  assign _03479_ = _03478_ | _03475_;
  assign _03480_ = _03479_ | _03472_;
  assign _03481_ = sel_oi_one_hot_i[136] & i[132];
  assign _03482_ = sel_oi_one_hot_i[137] & i[148];
  assign _03483_ = _03482_ | _03481_;
  assign _03484_ = sel_oi_one_hot_i[138] & i[164];
  assign _03485_ = sel_oi_one_hot_i[139] & i[180];
  assign _03486_ = _03485_ | _03484_;
  assign _03487_ = _03486_ | _03483_;
  assign _03488_ = sel_oi_one_hot_i[140] & i[196];
  assign _03489_ = sel_oi_one_hot_i[141] & i[212];
  assign _03490_ = _03489_ | _03488_;
  assign _03491_ = sel_oi_one_hot_i[142] & i[228];
  assign _03492_ = sel_oi_one_hot_i[143] & i[244];
  assign _03493_ = _03492_ | _03491_;
  assign _03494_ = _03493_ | _03490_;
  assign _03495_ = _03494_ | _03487_;
  assign o[132] = _03495_ | _03480_;
  assign _03496_ = sel_oi_one_hot_i[128] & i[3];
  assign _03497_ = sel_oi_one_hot_i[129] & i[19];
  assign _03498_ = _03497_ | _03496_;
  assign _03499_ = sel_oi_one_hot_i[130] & i[35];
  assign _03500_ = sel_oi_one_hot_i[131] & i[51];
  assign _03501_ = _03500_ | _03499_;
  assign _03502_ = _03501_ | _03498_;
  assign _03503_ = sel_oi_one_hot_i[132] & i[67];
  assign _03504_ = sel_oi_one_hot_i[133] & i[83];
  assign _03505_ = _03504_ | _03503_;
  assign _03506_ = sel_oi_one_hot_i[134] & i[99];
  assign _03507_ = sel_oi_one_hot_i[135] & i[115];
  assign _03508_ = _03507_ | _03506_;
  assign _03509_ = _03508_ | _03505_;
  assign _03510_ = _03509_ | _03502_;
  assign _03511_ = sel_oi_one_hot_i[136] & i[131];
  assign _03512_ = sel_oi_one_hot_i[137] & i[147];
  assign _03513_ = _03512_ | _03511_;
  assign _03514_ = sel_oi_one_hot_i[138] & i[163];
  assign _03515_ = sel_oi_one_hot_i[139] & i[179];
  assign _03516_ = _03515_ | _03514_;
  assign _03517_ = _03516_ | _03513_;
  assign _03518_ = sel_oi_one_hot_i[140] & i[195];
  assign _03519_ = sel_oi_one_hot_i[141] & i[211];
  assign _03520_ = _03519_ | _03518_;
  assign _03521_ = sel_oi_one_hot_i[142] & i[227];
  assign _03522_ = sel_oi_one_hot_i[143] & i[243];
  assign _03523_ = _03522_ | _03521_;
  assign _03524_ = _03523_ | _03520_;
  assign _03525_ = _03524_ | _03517_;
  assign o[131] = _03525_ | _03510_;
  assign _03526_ = sel_oi_one_hot_i[128] & i[2];
  assign _03527_ = sel_oi_one_hot_i[129] & i[18];
  assign _03528_ = _03527_ | _03526_;
  assign _03529_ = sel_oi_one_hot_i[130] & i[34];
  assign _03530_ = sel_oi_one_hot_i[131] & i[50];
  assign _03531_ = _03530_ | _03529_;
  assign _03532_ = _03531_ | _03528_;
  assign _03533_ = sel_oi_one_hot_i[132] & i[66];
  assign _03534_ = sel_oi_one_hot_i[133] & i[82];
  assign _03535_ = _03534_ | _03533_;
  assign _03536_ = sel_oi_one_hot_i[134] & i[98];
  assign _03537_ = sel_oi_one_hot_i[135] & i[114];
  assign _03538_ = _03537_ | _03536_;
  assign _03539_ = _03538_ | _03535_;
  assign _03540_ = _03539_ | _03532_;
  assign _03541_ = sel_oi_one_hot_i[136] & i[130];
  assign _03542_ = sel_oi_one_hot_i[137] & i[146];
  assign _03543_ = _03542_ | _03541_;
  assign _03544_ = sel_oi_one_hot_i[138] & i[162];
  assign _03545_ = sel_oi_one_hot_i[139] & i[178];
  assign _03546_ = _03545_ | _03544_;
  assign _03547_ = _03546_ | _03543_;
  assign _03548_ = sel_oi_one_hot_i[140] & i[194];
  assign _03549_ = sel_oi_one_hot_i[141] & i[210];
  assign _03550_ = _03549_ | _03548_;
  assign _03551_ = sel_oi_one_hot_i[142] & i[226];
  assign _03552_ = sel_oi_one_hot_i[143] & i[242];
  assign _03553_ = _03552_ | _03551_;
  assign _03554_ = _03553_ | _03550_;
  assign _03555_ = _03554_ | _03547_;
  assign o[130] = _03555_ | _03540_;
  assign _03556_ = sel_oi_one_hot_i[128] & i[1];
  assign _03557_ = sel_oi_one_hot_i[129] & i[17];
  assign _03558_ = _03557_ | _03556_;
  assign _03559_ = sel_oi_one_hot_i[130] & i[33];
  assign _03560_ = sel_oi_one_hot_i[131] & i[49];
  assign _03561_ = _03560_ | _03559_;
  assign _03562_ = _03561_ | _03558_;
  assign _03563_ = sel_oi_one_hot_i[132] & i[65];
  assign _03564_ = sel_oi_one_hot_i[133] & i[81];
  assign _03565_ = _03564_ | _03563_;
  assign _03566_ = sel_oi_one_hot_i[134] & i[97];
  assign _03567_ = sel_oi_one_hot_i[135] & i[113];
  assign _03568_ = _03567_ | _03566_;
  assign _03569_ = _03568_ | _03565_;
  assign _03570_ = _03569_ | _03562_;
  assign _03571_ = sel_oi_one_hot_i[136] & i[129];
  assign _03572_ = sel_oi_one_hot_i[137] & i[145];
  assign _03573_ = _03572_ | _03571_;
  assign _03574_ = sel_oi_one_hot_i[138] & i[161];
  assign _03575_ = sel_oi_one_hot_i[139] & i[177];
  assign _03576_ = _03575_ | _03574_;
  assign _03577_ = _03576_ | _03573_;
  assign _03578_ = sel_oi_one_hot_i[140] & i[193];
  assign _03579_ = sel_oi_one_hot_i[141] & i[209];
  assign _03580_ = _03579_ | _03578_;
  assign _03581_ = sel_oi_one_hot_i[142] & i[225];
  assign _03582_ = sel_oi_one_hot_i[143] & i[241];
  assign _03583_ = _03582_ | _03581_;
  assign _03584_ = _03583_ | _03580_;
  assign _03585_ = _03584_ | _03577_;
  assign o[129] = _03585_ | _03570_;
  assign _03586_ = sel_oi_one_hot_i[128] & i[0];
  assign _03587_ = sel_oi_one_hot_i[129] & i[16];
  assign _03588_ = _03587_ | _03586_;
  assign _03589_ = sel_oi_one_hot_i[130] & i[32];
  assign _03590_ = sel_oi_one_hot_i[131] & i[48];
  assign _03591_ = _03590_ | _03589_;
  assign _03592_ = _03591_ | _03588_;
  assign _03593_ = sel_oi_one_hot_i[132] & i[64];
  assign _03594_ = sel_oi_one_hot_i[133] & i[80];
  assign _03595_ = _03594_ | _03593_;
  assign _03596_ = sel_oi_one_hot_i[134] & i[96];
  assign _03597_ = sel_oi_one_hot_i[135] & i[112];
  assign _03598_ = _03597_ | _03596_;
  assign _03599_ = _03598_ | _03595_;
  assign _03600_ = _03599_ | _03592_;
  assign _03601_ = sel_oi_one_hot_i[136] & i[128];
  assign _03602_ = sel_oi_one_hot_i[137] & i[144];
  assign _03603_ = _03602_ | _03601_;
  assign _03604_ = sel_oi_one_hot_i[138] & i[160];
  assign _03605_ = sel_oi_one_hot_i[139] & i[176];
  assign _03606_ = _03605_ | _03604_;
  assign _03607_ = _03606_ | _03603_;
  assign _03608_ = sel_oi_one_hot_i[140] & i[192];
  assign _03609_ = sel_oi_one_hot_i[141] & i[208];
  assign _03610_ = _03609_ | _03608_;
  assign _03611_ = sel_oi_one_hot_i[142] & i[224];
  assign _03612_ = sel_oi_one_hot_i[143] & i[240];
  assign _03613_ = _03612_ | _03611_;
  assign _03614_ = _03613_ | _03610_;
  assign _03615_ = _03614_ | _03607_;
  assign o[128] = _03615_ | _03600_;
  assign _03616_ = sel_oi_one_hot_i[144] & i[15];
  assign _03617_ = sel_oi_one_hot_i[145] & i[31];
  assign _03618_ = _03617_ | _03616_;
  assign _03619_ = sel_oi_one_hot_i[146] & i[47];
  assign _03620_ = sel_oi_one_hot_i[147] & i[63];
  assign _03621_ = _03620_ | _03619_;
  assign _03622_ = _03621_ | _03618_;
  assign _03623_ = sel_oi_one_hot_i[148] & i[79];
  assign _03624_ = sel_oi_one_hot_i[149] & i[95];
  assign _03625_ = _03624_ | _03623_;
  assign _03626_ = sel_oi_one_hot_i[150] & i[111];
  assign _03627_ = sel_oi_one_hot_i[151] & i[127];
  assign _03628_ = _03627_ | _03626_;
  assign _03629_ = _03628_ | _03625_;
  assign _03630_ = _03629_ | _03622_;
  assign _03631_ = sel_oi_one_hot_i[152] & i[143];
  assign _03632_ = sel_oi_one_hot_i[153] & i[159];
  assign _03633_ = _03632_ | _03631_;
  assign _03634_ = sel_oi_one_hot_i[154] & i[175];
  assign _03635_ = sel_oi_one_hot_i[155] & i[191];
  assign _03636_ = _03635_ | _03634_;
  assign _03637_ = _03636_ | _03633_;
  assign _03638_ = sel_oi_one_hot_i[156] & i[207];
  assign _03639_ = sel_oi_one_hot_i[157] & i[223];
  assign _03640_ = _03639_ | _03638_;
  assign _03641_ = sel_oi_one_hot_i[158] & i[239];
  assign _03642_ = sel_oi_one_hot_i[159] & i[255];
  assign _03643_ = _03642_ | _03641_;
  assign _03644_ = _03643_ | _03640_;
  assign _03645_ = _03644_ | _03637_;
  assign o[159] = _03645_ | _03630_;
  assign _03646_ = sel_oi_one_hot_i[144] & i[14];
  assign _03647_ = sel_oi_one_hot_i[145] & i[30];
  assign _03648_ = _03647_ | _03646_;
  assign _03649_ = sel_oi_one_hot_i[146] & i[46];
  assign _03650_ = sel_oi_one_hot_i[147] & i[62];
  assign _03651_ = _03650_ | _03649_;
  assign _03652_ = _03651_ | _03648_;
  assign _03653_ = sel_oi_one_hot_i[148] & i[78];
  assign _03654_ = sel_oi_one_hot_i[149] & i[94];
  assign _03655_ = _03654_ | _03653_;
  assign _03656_ = sel_oi_one_hot_i[150] & i[110];
  assign _03657_ = sel_oi_one_hot_i[151] & i[126];
  assign _03658_ = _03657_ | _03656_;
  assign _03659_ = _03658_ | _03655_;
  assign _03660_ = _03659_ | _03652_;
  assign _03661_ = sel_oi_one_hot_i[152] & i[142];
  assign _03662_ = sel_oi_one_hot_i[153] & i[158];
  assign _03663_ = _03662_ | _03661_;
  assign _03664_ = sel_oi_one_hot_i[154] & i[174];
  assign _03665_ = sel_oi_one_hot_i[155] & i[190];
  assign _03666_ = _03665_ | _03664_;
  assign _03667_ = _03666_ | _03663_;
  assign _03668_ = sel_oi_one_hot_i[156] & i[206];
  assign _03669_ = sel_oi_one_hot_i[157] & i[222];
  assign _03670_ = _03669_ | _03668_;
  assign _03671_ = sel_oi_one_hot_i[158] & i[238];
  assign _03672_ = sel_oi_one_hot_i[159] & i[254];
  assign _03673_ = _03672_ | _03671_;
  assign _03674_ = _03673_ | _03670_;
  assign _03675_ = _03674_ | _03667_;
  assign o[158] = _03675_ | _03660_;
  assign _03676_ = sel_oi_one_hot_i[144] & i[13];
  assign _03677_ = sel_oi_one_hot_i[145] & i[29];
  assign _03678_ = _03677_ | _03676_;
  assign _03679_ = sel_oi_one_hot_i[146] & i[45];
  assign _03680_ = sel_oi_one_hot_i[147] & i[61];
  assign _03681_ = _03680_ | _03679_;
  assign _03682_ = _03681_ | _03678_;
  assign _03683_ = sel_oi_one_hot_i[148] & i[77];
  assign _03684_ = sel_oi_one_hot_i[149] & i[93];
  assign _03685_ = _03684_ | _03683_;
  assign _03686_ = sel_oi_one_hot_i[150] & i[109];
  assign _03687_ = sel_oi_one_hot_i[151] & i[125];
  assign _03688_ = _03687_ | _03686_;
  assign _03689_ = _03688_ | _03685_;
  assign _03690_ = _03689_ | _03682_;
  assign _03691_ = sel_oi_one_hot_i[152] & i[141];
  assign _03692_ = sel_oi_one_hot_i[153] & i[157];
  assign _03693_ = _03692_ | _03691_;
  assign _03694_ = sel_oi_one_hot_i[154] & i[173];
  assign _03695_ = sel_oi_one_hot_i[155] & i[189];
  assign _03696_ = _03695_ | _03694_;
  assign _03697_ = _03696_ | _03693_;
  assign _03698_ = sel_oi_one_hot_i[156] & i[205];
  assign _03699_ = sel_oi_one_hot_i[157] & i[221];
  assign _03700_ = _03699_ | _03698_;
  assign _03701_ = sel_oi_one_hot_i[158] & i[237];
  assign _03702_ = sel_oi_one_hot_i[159] & i[253];
  assign _03703_ = _03702_ | _03701_;
  assign _03704_ = _03703_ | _03700_;
  assign _03705_ = _03704_ | _03697_;
  assign o[157] = _03705_ | _03690_;
  assign _03706_ = sel_oi_one_hot_i[144] & i[12];
  assign _03707_ = sel_oi_one_hot_i[145] & i[28];
  assign _03708_ = _03707_ | _03706_;
  assign _03709_ = sel_oi_one_hot_i[146] & i[44];
  assign _03710_ = sel_oi_one_hot_i[147] & i[60];
  assign _03711_ = _03710_ | _03709_;
  assign _03712_ = _03711_ | _03708_;
  assign _03713_ = sel_oi_one_hot_i[148] & i[76];
  assign _03714_ = sel_oi_one_hot_i[149] & i[92];
  assign _03715_ = _03714_ | _03713_;
  assign _03716_ = sel_oi_one_hot_i[150] & i[108];
  assign _03717_ = sel_oi_one_hot_i[151] & i[124];
  assign _03718_ = _03717_ | _03716_;
  assign _03719_ = _03718_ | _03715_;
  assign _03720_ = _03719_ | _03712_;
  assign _03721_ = sel_oi_one_hot_i[152] & i[140];
  assign _03722_ = sel_oi_one_hot_i[153] & i[156];
  assign _03723_ = _03722_ | _03721_;
  assign _03724_ = sel_oi_one_hot_i[154] & i[172];
  assign _03725_ = sel_oi_one_hot_i[155] & i[188];
  assign _03726_ = _03725_ | _03724_;
  assign _03727_ = _03726_ | _03723_;
  assign _03728_ = sel_oi_one_hot_i[156] & i[204];
  assign _03729_ = sel_oi_one_hot_i[157] & i[220];
  assign _03730_ = _03729_ | _03728_;
  assign _03731_ = sel_oi_one_hot_i[158] & i[236];
  assign _03732_ = sel_oi_one_hot_i[159] & i[252];
  assign _03733_ = _03732_ | _03731_;
  assign _03734_ = _03733_ | _03730_;
  assign _03735_ = _03734_ | _03727_;
  assign o[156] = _03735_ | _03720_;
  assign _03736_ = sel_oi_one_hot_i[144] & i[11];
  assign _03737_ = sel_oi_one_hot_i[145] & i[27];
  assign _03738_ = _03737_ | _03736_;
  assign _03739_ = sel_oi_one_hot_i[146] & i[43];
  assign _03740_ = sel_oi_one_hot_i[147] & i[59];
  assign _03741_ = _03740_ | _03739_;
  assign _03742_ = _03741_ | _03738_;
  assign _03743_ = sel_oi_one_hot_i[148] & i[75];
  assign _03744_ = sel_oi_one_hot_i[149] & i[91];
  assign _03745_ = _03744_ | _03743_;
  assign _03746_ = sel_oi_one_hot_i[150] & i[107];
  assign _03747_ = sel_oi_one_hot_i[151] & i[123];
  assign _03748_ = _03747_ | _03746_;
  assign _03749_ = _03748_ | _03745_;
  assign _03750_ = _03749_ | _03742_;
  assign _03751_ = sel_oi_one_hot_i[152] & i[139];
  assign _03752_ = sel_oi_one_hot_i[153] & i[155];
  assign _03753_ = _03752_ | _03751_;
  assign _03754_ = sel_oi_one_hot_i[154] & i[171];
  assign _03755_ = sel_oi_one_hot_i[155] & i[187];
  assign _03756_ = _03755_ | _03754_;
  assign _03757_ = _03756_ | _03753_;
  assign _03758_ = sel_oi_one_hot_i[156] & i[203];
  assign _03759_ = sel_oi_one_hot_i[157] & i[219];
  assign _03760_ = _03759_ | _03758_;
  assign _03761_ = sel_oi_one_hot_i[158] & i[235];
  assign _03762_ = sel_oi_one_hot_i[159] & i[251];
  assign _03763_ = _03762_ | _03761_;
  assign _03764_ = _03763_ | _03760_;
  assign _03765_ = _03764_ | _03757_;
  assign o[155] = _03765_ | _03750_;
  assign _03766_ = sel_oi_one_hot_i[144] & i[10];
  assign _03767_ = sel_oi_one_hot_i[145] & i[26];
  assign _03768_ = _03767_ | _03766_;
  assign _03769_ = sel_oi_one_hot_i[146] & i[42];
  assign _03770_ = sel_oi_one_hot_i[147] & i[58];
  assign _03771_ = _03770_ | _03769_;
  assign _03772_ = _03771_ | _03768_;
  assign _03773_ = sel_oi_one_hot_i[148] & i[74];
  assign _03774_ = sel_oi_one_hot_i[149] & i[90];
  assign _03775_ = _03774_ | _03773_;
  assign _03776_ = sel_oi_one_hot_i[150] & i[106];
  assign _03777_ = sel_oi_one_hot_i[151] & i[122];
  assign _03778_ = _03777_ | _03776_;
  assign _03779_ = _03778_ | _03775_;
  assign _03780_ = _03779_ | _03772_;
  assign _03781_ = sel_oi_one_hot_i[152] & i[138];
  assign _03782_ = sel_oi_one_hot_i[153] & i[154];
  assign _03783_ = _03782_ | _03781_;
  assign _03784_ = sel_oi_one_hot_i[154] & i[170];
  assign _03785_ = sel_oi_one_hot_i[155] & i[186];
  assign _03786_ = _03785_ | _03784_;
  assign _03787_ = _03786_ | _03783_;
  assign _03788_ = sel_oi_one_hot_i[156] & i[202];
  assign _03789_ = sel_oi_one_hot_i[157] & i[218];
  assign _03790_ = _03789_ | _03788_;
  assign _03791_ = sel_oi_one_hot_i[158] & i[234];
  assign _03792_ = sel_oi_one_hot_i[159] & i[250];
  assign _03793_ = _03792_ | _03791_;
  assign _03794_ = _03793_ | _03790_;
  assign _03795_ = _03794_ | _03787_;
  assign o[154] = _03795_ | _03780_;
  assign _03796_ = sel_oi_one_hot_i[144] & i[9];
  assign _03797_ = sel_oi_one_hot_i[145] & i[25];
  assign _03798_ = _03797_ | _03796_;
  assign _03799_ = sel_oi_one_hot_i[146] & i[41];
  assign _03800_ = sel_oi_one_hot_i[147] & i[57];
  assign _03801_ = _03800_ | _03799_;
  assign _03802_ = _03801_ | _03798_;
  assign _03803_ = sel_oi_one_hot_i[148] & i[73];
  assign _03804_ = sel_oi_one_hot_i[149] & i[89];
  assign _03805_ = _03804_ | _03803_;
  assign _03806_ = sel_oi_one_hot_i[150] & i[105];
  assign _03807_ = sel_oi_one_hot_i[151] & i[121];
  assign _03808_ = _03807_ | _03806_;
  assign _03809_ = _03808_ | _03805_;
  assign _03810_ = _03809_ | _03802_;
  assign _03811_ = sel_oi_one_hot_i[152] & i[137];
  assign _03812_ = sel_oi_one_hot_i[153] & i[153];
  assign _03813_ = _03812_ | _03811_;
  assign _03814_ = sel_oi_one_hot_i[154] & i[169];
  assign _03815_ = sel_oi_one_hot_i[155] & i[185];
  assign _03816_ = _03815_ | _03814_;
  assign _03817_ = _03816_ | _03813_;
  assign _03818_ = sel_oi_one_hot_i[156] & i[201];
  assign _03819_ = sel_oi_one_hot_i[157] & i[217];
  assign _03820_ = _03819_ | _03818_;
  assign _03821_ = sel_oi_one_hot_i[158] & i[233];
  assign _03822_ = sel_oi_one_hot_i[159] & i[249];
  assign _03823_ = _03822_ | _03821_;
  assign _03824_ = _03823_ | _03820_;
  assign _03825_ = _03824_ | _03817_;
  assign o[153] = _03825_ | _03810_;
  assign _03826_ = sel_oi_one_hot_i[144] & i[8];
  assign _03827_ = sel_oi_one_hot_i[145] & i[24];
  assign _03828_ = _03827_ | _03826_;
  assign _03829_ = sel_oi_one_hot_i[146] & i[40];
  assign _03830_ = sel_oi_one_hot_i[147] & i[56];
  assign _03831_ = _03830_ | _03829_;
  assign _03832_ = _03831_ | _03828_;
  assign _03833_ = sel_oi_one_hot_i[148] & i[72];
  assign _03834_ = sel_oi_one_hot_i[149] & i[88];
  assign _03835_ = _03834_ | _03833_;
  assign _03836_ = sel_oi_one_hot_i[150] & i[104];
  assign _03837_ = sel_oi_one_hot_i[151] & i[120];
  assign _03838_ = _03837_ | _03836_;
  assign _03839_ = _03838_ | _03835_;
  assign _03840_ = _03839_ | _03832_;
  assign _03841_ = sel_oi_one_hot_i[152] & i[136];
  assign _03842_ = sel_oi_one_hot_i[153] & i[152];
  assign _03843_ = _03842_ | _03841_;
  assign _03844_ = sel_oi_one_hot_i[154] & i[168];
  assign _03845_ = sel_oi_one_hot_i[155] & i[184];
  assign _03846_ = _03845_ | _03844_;
  assign _03847_ = _03846_ | _03843_;
  assign _03848_ = sel_oi_one_hot_i[156] & i[200];
  assign _03849_ = sel_oi_one_hot_i[157] & i[216];
  assign _03850_ = _03849_ | _03848_;
  assign _03851_ = sel_oi_one_hot_i[158] & i[232];
  assign _03852_ = sel_oi_one_hot_i[159] & i[248];
  assign _03853_ = _03852_ | _03851_;
  assign _03854_ = _03853_ | _03850_;
  assign _03855_ = _03854_ | _03847_;
  assign o[152] = _03855_ | _03840_;
  assign _03856_ = sel_oi_one_hot_i[144] & i[7];
  assign _03857_ = sel_oi_one_hot_i[145] & i[23];
  assign _03858_ = _03857_ | _03856_;
  assign _03859_ = sel_oi_one_hot_i[146] & i[39];
  assign _03860_ = sel_oi_one_hot_i[147] & i[55];
  assign _03861_ = _03860_ | _03859_;
  assign _03862_ = _03861_ | _03858_;
  assign _03863_ = sel_oi_one_hot_i[148] & i[71];
  assign _03864_ = sel_oi_one_hot_i[149] & i[87];
  assign _03865_ = _03864_ | _03863_;
  assign _03866_ = sel_oi_one_hot_i[150] & i[103];
  assign _03867_ = sel_oi_one_hot_i[151] & i[119];
  assign _03868_ = _03867_ | _03866_;
  assign _03869_ = _03868_ | _03865_;
  assign _03870_ = _03869_ | _03862_;
  assign _03871_ = sel_oi_one_hot_i[152] & i[135];
  assign _03872_ = sel_oi_one_hot_i[153] & i[151];
  assign _03873_ = _03872_ | _03871_;
  assign _03874_ = sel_oi_one_hot_i[154] & i[167];
  assign _03875_ = sel_oi_one_hot_i[155] & i[183];
  assign _03876_ = _03875_ | _03874_;
  assign _03877_ = _03876_ | _03873_;
  assign _03878_ = sel_oi_one_hot_i[156] & i[199];
  assign _03879_ = sel_oi_one_hot_i[157] & i[215];
  assign _03880_ = _03879_ | _03878_;
  assign _03881_ = sel_oi_one_hot_i[158] & i[231];
  assign _03882_ = sel_oi_one_hot_i[159] & i[247];
  assign _03883_ = _03882_ | _03881_;
  assign _03884_ = _03883_ | _03880_;
  assign _03885_ = _03884_ | _03877_;
  assign o[151] = _03885_ | _03870_;
  assign _03886_ = sel_oi_one_hot_i[144] & i[6];
  assign _03887_ = sel_oi_one_hot_i[145] & i[22];
  assign _03888_ = _03887_ | _03886_;
  assign _03889_ = sel_oi_one_hot_i[146] & i[38];
  assign _03890_ = sel_oi_one_hot_i[147] & i[54];
  assign _03891_ = _03890_ | _03889_;
  assign _03892_ = _03891_ | _03888_;
  assign _03893_ = sel_oi_one_hot_i[148] & i[70];
  assign _03894_ = sel_oi_one_hot_i[149] & i[86];
  assign _03895_ = _03894_ | _03893_;
  assign _03896_ = sel_oi_one_hot_i[150] & i[102];
  assign _03897_ = sel_oi_one_hot_i[151] & i[118];
  assign _03898_ = _03897_ | _03896_;
  assign _03899_ = _03898_ | _03895_;
  assign _03900_ = _03899_ | _03892_;
  assign _03901_ = sel_oi_one_hot_i[152] & i[134];
  assign _03902_ = sel_oi_one_hot_i[153] & i[150];
  assign _03903_ = _03902_ | _03901_;
  assign _03904_ = sel_oi_one_hot_i[154] & i[166];
  assign _03905_ = sel_oi_one_hot_i[155] & i[182];
  assign _03906_ = _03905_ | _03904_;
  assign _03907_ = _03906_ | _03903_;
  assign _03908_ = sel_oi_one_hot_i[156] & i[198];
  assign _03909_ = sel_oi_one_hot_i[157] & i[214];
  assign _03910_ = _03909_ | _03908_;
  assign _03911_ = sel_oi_one_hot_i[158] & i[230];
  assign _03912_ = sel_oi_one_hot_i[159] & i[246];
  assign _03913_ = _03912_ | _03911_;
  assign _03914_ = _03913_ | _03910_;
  assign _03915_ = _03914_ | _03907_;
  assign o[150] = _03915_ | _03900_;
  assign _03916_ = sel_oi_one_hot_i[144] & i[5];
  assign _03917_ = sel_oi_one_hot_i[145] & i[21];
  assign _03918_ = _03917_ | _03916_;
  assign _03919_ = sel_oi_one_hot_i[146] & i[37];
  assign _03920_ = sel_oi_one_hot_i[147] & i[53];
  assign _03921_ = _03920_ | _03919_;
  assign _03922_ = _03921_ | _03918_;
  assign _03923_ = sel_oi_one_hot_i[148] & i[69];
  assign _03924_ = sel_oi_one_hot_i[149] & i[85];
  assign _03925_ = _03924_ | _03923_;
  assign _03926_ = sel_oi_one_hot_i[150] & i[101];
  assign _03927_ = sel_oi_one_hot_i[151] & i[117];
  assign _03928_ = _03927_ | _03926_;
  assign _03929_ = _03928_ | _03925_;
  assign _03930_ = _03929_ | _03922_;
  assign _03931_ = sel_oi_one_hot_i[152] & i[133];
  assign _03932_ = sel_oi_one_hot_i[153] & i[149];
  assign _03933_ = _03932_ | _03931_;
  assign _03934_ = sel_oi_one_hot_i[154] & i[165];
  assign _03935_ = sel_oi_one_hot_i[155] & i[181];
  assign _03936_ = _03935_ | _03934_;
  assign _03937_ = _03936_ | _03933_;
  assign _03938_ = sel_oi_one_hot_i[156] & i[197];
  assign _03939_ = sel_oi_one_hot_i[157] & i[213];
  assign _03940_ = _03939_ | _03938_;
  assign _03941_ = sel_oi_one_hot_i[158] & i[229];
  assign _03942_ = sel_oi_one_hot_i[159] & i[245];
  assign _03943_ = _03942_ | _03941_;
  assign _03944_ = _03943_ | _03940_;
  assign _03945_ = _03944_ | _03937_;
  assign o[149] = _03945_ | _03930_;
  assign _03946_ = sel_oi_one_hot_i[144] & i[4];
  assign _03947_ = sel_oi_one_hot_i[145] & i[20];
  assign _03948_ = _03947_ | _03946_;
  assign _03949_ = sel_oi_one_hot_i[146] & i[36];
  assign _03950_ = sel_oi_one_hot_i[147] & i[52];
  assign _03951_ = _03950_ | _03949_;
  assign _03952_ = _03951_ | _03948_;
  assign _03953_ = sel_oi_one_hot_i[148] & i[68];
  assign _03954_ = sel_oi_one_hot_i[149] & i[84];
  assign _03955_ = _03954_ | _03953_;
  assign _03956_ = sel_oi_one_hot_i[150] & i[100];
  assign _03957_ = sel_oi_one_hot_i[151] & i[116];
  assign _03958_ = _03957_ | _03956_;
  assign _03959_ = _03958_ | _03955_;
  assign _03960_ = _03959_ | _03952_;
  assign _03961_ = sel_oi_one_hot_i[152] & i[132];
  assign _03962_ = sel_oi_one_hot_i[153] & i[148];
  assign _03963_ = _03962_ | _03961_;
  assign _03964_ = sel_oi_one_hot_i[154] & i[164];
  assign _03965_ = sel_oi_one_hot_i[155] & i[180];
  assign _03966_ = _03965_ | _03964_;
  assign _03967_ = _03966_ | _03963_;
  assign _03968_ = sel_oi_one_hot_i[156] & i[196];
  assign _03969_ = sel_oi_one_hot_i[157] & i[212];
  assign _03970_ = _03969_ | _03968_;
  assign _03971_ = sel_oi_one_hot_i[158] & i[228];
  assign _03972_ = sel_oi_one_hot_i[159] & i[244];
  assign _03973_ = _03972_ | _03971_;
  assign _03974_ = _03973_ | _03970_;
  assign _03975_ = _03974_ | _03967_;
  assign o[148] = _03975_ | _03960_;
  assign _03976_ = sel_oi_one_hot_i[144] & i[3];
  assign _03977_ = sel_oi_one_hot_i[145] & i[19];
  assign _03978_ = _03977_ | _03976_;
  assign _03979_ = sel_oi_one_hot_i[146] & i[35];
  assign _03980_ = sel_oi_one_hot_i[147] & i[51];
  assign _03981_ = _03980_ | _03979_;
  assign _03982_ = _03981_ | _03978_;
  assign _03983_ = sel_oi_one_hot_i[148] & i[67];
  assign _03984_ = sel_oi_one_hot_i[149] & i[83];
  assign _03985_ = _03984_ | _03983_;
  assign _03986_ = sel_oi_one_hot_i[150] & i[99];
  assign _03987_ = sel_oi_one_hot_i[151] & i[115];
  assign _03988_ = _03987_ | _03986_;
  assign _03989_ = _03988_ | _03985_;
  assign _03990_ = _03989_ | _03982_;
  assign _03991_ = sel_oi_one_hot_i[152] & i[131];
  assign _03992_ = sel_oi_one_hot_i[153] & i[147];
  assign _03993_ = _03992_ | _03991_;
  assign _03994_ = sel_oi_one_hot_i[154] & i[163];
  assign _03995_ = sel_oi_one_hot_i[155] & i[179];
  assign _03996_ = _03995_ | _03994_;
  assign _03997_ = _03996_ | _03993_;
  assign _03998_ = sel_oi_one_hot_i[156] & i[195];
  assign _03999_ = sel_oi_one_hot_i[157] & i[211];
  assign _04000_ = _03999_ | _03998_;
  assign _04001_ = sel_oi_one_hot_i[158] & i[227];
  assign _04002_ = sel_oi_one_hot_i[159] & i[243];
  assign _04003_ = _04002_ | _04001_;
  assign _04004_ = _04003_ | _04000_;
  assign _04005_ = _04004_ | _03997_;
  assign o[147] = _04005_ | _03990_;
  assign _04006_ = sel_oi_one_hot_i[144] & i[2];
  assign _04007_ = sel_oi_one_hot_i[145] & i[18];
  assign _04008_ = _04007_ | _04006_;
  assign _04009_ = sel_oi_one_hot_i[146] & i[34];
  assign _04010_ = sel_oi_one_hot_i[147] & i[50];
  assign _04011_ = _04010_ | _04009_;
  assign _04012_ = _04011_ | _04008_;
  assign _04013_ = sel_oi_one_hot_i[148] & i[66];
  assign _04014_ = sel_oi_one_hot_i[149] & i[82];
  assign _04015_ = _04014_ | _04013_;
  assign _04016_ = sel_oi_one_hot_i[150] & i[98];
  assign _04017_ = sel_oi_one_hot_i[151] & i[114];
  assign _04018_ = _04017_ | _04016_;
  assign _04019_ = _04018_ | _04015_;
  assign _04020_ = _04019_ | _04012_;
  assign _04021_ = sel_oi_one_hot_i[152] & i[130];
  assign _04022_ = sel_oi_one_hot_i[153] & i[146];
  assign _04023_ = _04022_ | _04021_;
  assign _04024_ = sel_oi_one_hot_i[154] & i[162];
  assign _04025_ = sel_oi_one_hot_i[155] & i[178];
  assign _04026_ = _04025_ | _04024_;
  assign _04027_ = _04026_ | _04023_;
  assign _04028_ = sel_oi_one_hot_i[156] & i[194];
  assign _04029_ = sel_oi_one_hot_i[157] & i[210];
  assign _04030_ = _04029_ | _04028_;
  assign _04031_ = sel_oi_one_hot_i[158] & i[226];
  assign _04032_ = sel_oi_one_hot_i[159] & i[242];
  assign _04033_ = _04032_ | _04031_;
  assign _04034_ = _04033_ | _04030_;
  assign _04035_ = _04034_ | _04027_;
  assign o[146] = _04035_ | _04020_;
  assign _04036_ = sel_oi_one_hot_i[144] & i[1];
  assign _04037_ = sel_oi_one_hot_i[145] & i[17];
  assign _04038_ = _04037_ | _04036_;
  assign _04039_ = sel_oi_one_hot_i[146] & i[33];
  assign _04040_ = sel_oi_one_hot_i[147] & i[49];
  assign _04041_ = _04040_ | _04039_;
  assign _04042_ = _04041_ | _04038_;
  assign _04043_ = sel_oi_one_hot_i[148] & i[65];
  assign _04044_ = sel_oi_one_hot_i[149] & i[81];
  assign _04045_ = _04044_ | _04043_;
  assign _04046_ = sel_oi_one_hot_i[150] & i[97];
  assign _04047_ = sel_oi_one_hot_i[151] & i[113];
  assign _04048_ = _04047_ | _04046_;
  assign _04049_ = _04048_ | _04045_;
  assign _04050_ = _04049_ | _04042_;
  assign _04051_ = sel_oi_one_hot_i[152] & i[129];
  assign _04052_ = sel_oi_one_hot_i[153] & i[145];
  assign _04053_ = _04052_ | _04051_;
  assign _04054_ = sel_oi_one_hot_i[154] & i[161];
  assign _04055_ = sel_oi_one_hot_i[155] & i[177];
  assign _04056_ = _04055_ | _04054_;
  assign _04057_ = _04056_ | _04053_;
  assign _04058_ = sel_oi_one_hot_i[156] & i[193];
  assign _04059_ = sel_oi_one_hot_i[157] & i[209];
  assign _04060_ = _04059_ | _04058_;
  assign _04061_ = sel_oi_one_hot_i[158] & i[225];
  assign _04062_ = sel_oi_one_hot_i[159] & i[241];
  assign _04063_ = _04062_ | _04061_;
  assign _04064_ = _04063_ | _04060_;
  assign _04065_ = _04064_ | _04057_;
  assign o[145] = _04065_ | _04050_;
  assign _04066_ = sel_oi_one_hot_i[144] & i[0];
  assign _04067_ = sel_oi_one_hot_i[145] & i[16];
  assign _04068_ = _04067_ | _04066_;
  assign _04069_ = sel_oi_one_hot_i[146] & i[32];
  assign _04070_ = sel_oi_one_hot_i[147] & i[48];
  assign _04071_ = _04070_ | _04069_;
  assign _04072_ = _04071_ | _04068_;
  assign _04073_ = sel_oi_one_hot_i[148] & i[64];
  assign _04074_ = sel_oi_one_hot_i[149] & i[80];
  assign _04075_ = _04074_ | _04073_;
  assign _04076_ = sel_oi_one_hot_i[150] & i[96];
  assign _04077_ = sel_oi_one_hot_i[151] & i[112];
  assign _04078_ = _04077_ | _04076_;
  assign _04079_ = _04078_ | _04075_;
  assign _04080_ = _04079_ | _04072_;
  assign _04081_ = sel_oi_one_hot_i[152] & i[128];
  assign _04082_ = sel_oi_one_hot_i[153] & i[144];
  assign _04083_ = _04082_ | _04081_;
  assign _04084_ = sel_oi_one_hot_i[154] & i[160];
  assign _04085_ = sel_oi_one_hot_i[155] & i[176];
  assign _04086_ = _04085_ | _04084_;
  assign _04087_ = _04086_ | _04083_;
  assign _04088_ = sel_oi_one_hot_i[156] & i[192];
  assign _04089_ = sel_oi_one_hot_i[157] & i[208];
  assign _04090_ = _04089_ | _04088_;
  assign _04091_ = sel_oi_one_hot_i[158] & i[224];
  assign _04092_ = sel_oi_one_hot_i[159] & i[240];
  assign _04093_ = _04092_ | _04091_;
  assign _04094_ = _04093_ | _04090_;
  assign _04095_ = _04094_ | _04087_;
  assign o[144] = _04095_ | _04080_;
  assign _04096_ = sel_oi_one_hot_i[160] & i[15];
  assign _04097_ = sel_oi_one_hot_i[161] & i[31];
  assign _04098_ = _04097_ | _04096_;
  assign _04099_ = sel_oi_one_hot_i[162] & i[47];
  assign _04100_ = sel_oi_one_hot_i[163] & i[63];
  assign _04101_ = _04100_ | _04099_;
  assign _04102_ = _04101_ | _04098_;
  assign _04103_ = sel_oi_one_hot_i[164] & i[79];
  assign _04104_ = sel_oi_one_hot_i[165] & i[95];
  assign _04105_ = _04104_ | _04103_;
  assign _04106_ = sel_oi_one_hot_i[166] & i[111];
  assign _04107_ = sel_oi_one_hot_i[167] & i[127];
  assign _04108_ = _04107_ | _04106_;
  assign _04109_ = _04108_ | _04105_;
  assign _04110_ = _04109_ | _04102_;
  assign _04111_ = sel_oi_one_hot_i[168] & i[143];
  assign _04112_ = sel_oi_one_hot_i[169] & i[159];
  assign _04113_ = _04112_ | _04111_;
  assign _04114_ = sel_oi_one_hot_i[170] & i[175];
  assign _04115_ = sel_oi_one_hot_i[171] & i[191];
  assign _04116_ = _04115_ | _04114_;
  assign _04117_ = _04116_ | _04113_;
  assign _04118_ = sel_oi_one_hot_i[172] & i[207];
  assign _04119_ = sel_oi_one_hot_i[173] & i[223];
  assign _04120_ = _04119_ | _04118_;
  assign _04121_ = sel_oi_one_hot_i[174] & i[239];
  assign _04122_ = sel_oi_one_hot_i[175] & i[255];
  assign _04123_ = _04122_ | _04121_;
  assign _04124_ = _04123_ | _04120_;
  assign _04125_ = _04124_ | _04117_;
  assign o[175] = _04125_ | _04110_;
  assign _04126_ = sel_oi_one_hot_i[160] & i[14];
  assign _04127_ = sel_oi_one_hot_i[161] & i[30];
  assign _04128_ = _04127_ | _04126_;
  assign _04129_ = sel_oi_one_hot_i[162] & i[46];
  assign _04130_ = sel_oi_one_hot_i[163] & i[62];
  assign _04131_ = _04130_ | _04129_;
  assign _04132_ = _04131_ | _04128_;
  assign _04133_ = sel_oi_one_hot_i[164] & i[78];
  assign _04134_ = sel_oi_one_hot_i[165] & i[94];
  assign _04135_ = _04134_ | _04133_;
  assign _04136_ = sel_oi_one_hot_i[166] & i[110];
  assign _04137_ = sel_oi_one_hot_i[167] & i[126];
  assign _04138_ = _04137_ | _04136_;
  assign _04139_ = _04138_ | _04135_;
  assign _04140_ = _04139_ | _04132_;
  assign _04141_ = sel_oi_one_hot_i[168] & i[142];
  assign _04142_ = sel_oi_one_hot_i[169] & i[158];
  assign _04143_ = _04142_ | _04141_;
  assign _04144_ = sel_oi_one_hot_i[170] & i[174];
  assign _04145_ = sel_oi_one_hot_i[171] & i[190];
  assign _04146_ = _04145_ | _04144_;
  assign _04147_ = _04146_ | _04143_;
  assign _04148_ = sel_oi_one_hot_i[172] & i[206];
  assign _04149_ = sel_oi_one_hot_i[173] & i[222];
  assign _04150_ = _04149_ | _04148_;
  assign _04151_ = sel_oi_one_hot_i[174] & i[238];
  assign _04152_ = sel_oi_one_hot_i[175] & i[254];
  assign _04153_ = _04152_ | _04151_;
  assign _04154_ = _04153_ | _04150_;
  assign _04155_ = _04154_ | _04147_;
  assign o[174] = _04155_ | _04140_;
  assign _04156_ = sel_oi_one_hot_i[160] & i[13];
  assign _04157_ = sel_oi_one_hot_i[161] & i[29];
  assign _04158_ = _04157_ | _04156_;
  assign _04159_ = sel_oi_one_hot_i[162] & i[45];
  assign _04160_ = sel_oi_one_hot_i[163] & i[61];
  assign _04161_ = _04160_ | _04159_;
  assign _04162_ = _04161_ | _04158_;
  assign _04163_ = sel_oi_one_hot_i[164] & i[77];
  assign _04164_ = sel_oi_one_hot_i[165] & i[93];
  assign _04165_ = _04164_ | _04163_;
  assign _04166_ = sel_oi_one_hot_i[166] & i[109];
  assign _04167_ = sel_oi_one_hot_i[167] & i[125];
  assign _04168_ = _04167_ | _04166_;
  assign _04169_ = _04168_ | _04165_;
  assign _04170_ = _04169_ | _04162_;
  assign _04171_ = sel_oi_one_hot_i[168] & i[141];
  assign _04172_ = sel_oi_one_hot_i[169] & i[157];
  assign _04173_ = _04172_ | _04171_;
  assign _04174_ = sel_oi_one_hot_i[170] & i[173];
  assign _04175_ = sel_oi_one_hot_i[171] & i[189];
  assign _04176_ = _04175_ | _04174_;
  assign _04177_ = _04176_ | _04173_;
  assign _04178_ = sel_oi_one_hot_i[172] & i[205];
  assign _04179_ = sel_oi_one_hot_i[173] & i[221];
  assign _04180_ = _04179_ | _04178_;
  assign _04181_ = sel_oi_one_hot_i[174] & i[237];
  assign _04182_ = sel_oi_one_hot_i[175] & i[253];
  assign _04183_ = _04182_ | _04181_;
  assign _04184_ = _04183_ | _04180_;
  assign _04185_ = _04184_ | _04177_;
  assign o[173] = _04185_ | _04170_;
  assign _04186_ = sel_oi_one_hot_i[160] & i[12];
  assign _04187_ = sel_oi_one_hot_i[161] & i[28];
  assign _04188_ = _04187_ | _04186_;
  assign _04189_ = sel_oi_one_hot_i[162] & i[44];
  assign _04190_ = sel_oi_one_hot_i[163] & i[60];
  assign _04191_ = _04190_ | _04189_;
  assign _04192_ = _04191_ | _04188_;
  assign _04193_ = sel_oi_one_hot_i[164] & i[76];
  assign _04194_ = sel_oi_one_hot_i[165] & i[92];
  assign _04195_ = _04194_ | _04193_;
  assign _04196_ = sel_oi_one_hot_i[166] & i[108];
  assign _04197_ = sel_oi_one_hot_i[167] & i[124];
  assign _04198_ = _04197_ | _04196_;
  assign _04199_ = _04198_ | _04195_;
  assign _04200_ = _04199_ | _04192_;
  assign _04201_ = sel_oi_one_hot_i[168] & i[140];
  assign _04202_ = sel_oi_one_hot_i[169] & i[156];
  assign _04203_ = _04202_ | _04201_;
  assign _04204_ = sel_oi_one_hot_i[170] & i[172];
  assign _04205_ = sel_oi_one_hot_i[171] & i[188];
  assign _04206_ = _04205_ | _04204_;
  assign _04207_ = _04206_ | _04203_;
  assign _04208_ = sel_oi_one_hot_i[172] & i[204];
  assign _04209_ = sel_oi_one_hot_i[173] & i[220];
  assign _04210_ = _04209_ | _04208_;
  assign _04211_ = sel_oi_one_hot_i[174] & i[236];
  assign _04212_ = sel_oi_one_hot_i[175] & i[252];
  assign _04213_ = _04212_ | _04211_;
  assign _04214_ = _04213_ | _04210_;
  assign _04215_ = _04214_ | _04207_;
  assign o[172] = _04215_ | _04200_;
  assign _04216_ = sel_oi_one_hot_i[160] & i[11];
  assign _04217_ = sel_oi_one_hot_i[161] & i[27];
  assign _04218_ = _04217_ | _04216_;
  assign _04219_ = sel_oi_one_hot_i[162] & i[43];
  assign _04220_ = sel_oi_one_hot_i[163] & i[59];
  assign _04221_ = _04220_ | _04219_;
  assign _04222_ = _04221_ | _04218_;
  assign _04223_ = sel_oi_one_hot_i[164] & i[75];
  assign _04224_ = sel_oi_one_hot_i[165] & i[91];
  assign _04225_ = _04224_ | _04223_;
  assign _04226_ = sel_oi_one_hot_i[166] & i[107];
  assign _04227_ = sel_oi_one_hot_i[167] & i[123];
  assign _04228_ = _04227_ | _04226_;
  assign _04229_ = _04228_ | _04225_;
  assign _04230_ = _04229_ | _04222_;
  assign _04231_ = sel_oi_one_hot_i[168] & i[139];
  assign _04232_ = sel_oi_one_hot_i[169] & i[155];
  assign _04233_ = _04232_ | _04231_;
  assign _04234_ = sel_oi_one_hot_i[170] & i[171];
  assign _04235_ = sel_oi_one_hot_i[171] & i[187];
  assign _04236_ = _04235_ | _04234_;
  assign _04237_ = _04236_ | _04233_;
  assign _04238_ = sel_oi_one_hot_i[172] & i[203];
  assign _04239_ = sel_oi_one_hot_i[173] & i[219];
  assign _04240_ = _04239_ | _04238_;
  assign _04241_ = sel_oi_one_hot_i[174] & i[235];
  assign _04242_ = sel_oi_one_hot_i[175] & i[251];
  assign _04243_ = _04242_ | _04241_;
  assign _04244_ = _04243_ | _04240_;
  assign _04245_ = _04244_ | _04237_;
  assign o[171] = _04245_ | _04230_;
  assign _04246_ = sel_oi_one_hot_i[160] & i[10];
  assign _04247_ = sel_oi_one_hot_i[161] & i[26];
  assign _04248_ = _04247_ | _04246_;
  assign _04249_ = sel_oi_one_hot_i[162] & i[42];
  assign _04250_ = sel_oi_one_hot_i[163] & i[58];
  assign _04251_ = _04250_ | _04249_;
  assign _04252_ = _04251_ | _04248_;
  assign _04253_ = sel_oi_one_hot_i[164] & i[74];
  assign _04254_ = sel_oi_one_hot_i[165] & i[90];
  assign _04255_ = _04254_ | _04253_;
  assign _04256_ = sel_oi_one_hot_i[166] & i[106];
  assign _04257_ = sel_oi_one_hot_i[167] & i[122];
  assign _04258_ = _04257_ | _04256_;
  assign _04259_ = _04258_ | _04255_;
  assign _04260_ = _04259_ | _04252_;
  assign _04261_ = sel_oi_one_hot_i[168] & i[138];
  assign _04262_ = sel_oi_one_hot_i[169] & i[154];
  assign _04263_ = _04262_ | _04261_;
  assign _04264_ = sel_oi_one_hot_i[170] & i[170];
  assign _04265_ = sel_oi_one_hot_i[171] & i[186];
  assign _04266_ = _04265_ | _04264_;
  assign _04267_ = _04266_ | _04263_;
  assign _04268_ = sel_oi_one_hot_i[172] & i[202];
  assign _04269_ = sel_oi_one_hot_i[173] & i[218];
  assign _04270_ = _04269_ | _04268_;
  assign _04271_ = sel_oi_one_hot_i[174] & i[234];
  assign _04272_ = sel_oi_one_hot_i[175] & i[250];
  assign _04273_ = _04272_ | _04271_;
  assign _04274_ = _04273_ | _04270_;
  assign _04275_ = _04274_ | _04267_;
  assign o[170] = _04275_ | _04260_;
  assign _04276_ = sel_oi_one_hot_i[160] & i[9];
  assign _04277_ = sel_oi_one_hot_i[161] & i[25];
  assign _04278_ = _04277_ | _04276_;
  assign _04279_ = sel_oi_one_hot_i[162] & i[41];
  assign _04280_ = sel_oi_one_hot_i[163] & i[57];
  assign _04281_ = _04280_ | _04279_;
  assign _04282_ = _04281_ | _04278_;
  assign _04283_ = sel_oi_one_hot_i[164] & i[73];
  assign _04284_ = sel_oi_one_hot_i[165] & i[89];
  assign _04285_ = _04284_ | _04283_;
  assign _04286_ = sel_oi_one_hot_i[166] & i[105];
  assign _04287_ = sel_oi_one_hot_i[167] & i[121];
  assign _04288_ = _04287_ | _04286_;
  assign _04289_ = _04288_ | _04285_;
  assign _04290_ = _04289_ | _04282_;
  assign _04291_ = sel_oi_one_hot_i[168] & i[137];
  assign _04292_ = sel_oi_one_hot_i[169] & i[153];
  assign _04293_ = _04292_ | _04291_;
  assign _04294_ = sel_oi_one_hot_i[170] & i[169];
  assign _04295_ = sel_oi_one_hot_i[171] & i[185];
  assign _04296_ = _04295_ | _04294_;
  assign _04297_ = _04296_ | _04293_;
  assign _04298_ = sel_oi_one_hot_i[172] & i[201];
  assign _04299_ = sel_oi_one_hot_i[173] & i[217];
  assign _04300_ = _04299_ | _04298_;
  assign _04301_ = sel_oi_one_hot_i[174] & i[233];
  assign _04302_ = sel_oi_one_hot_i[175] & i[249];
  assign _04303_ = _04302_ | _04301_;
  assign _04304_ = _04303_ | _04300_;
  assign _04305_ = _04304_ | _04297_;
  assign o[169] = _04305_ | _04290_;
  assign _04306_ = sel_oi_one_hot_i[160] & i[8];
  assign _04307_ = sel_oi_one_hot_i[161] & i[24];
  assign _04308_ = _04307_ | _04306_;
  assign _04309_ = sel_oi_one_hot_i[162] & i[40];
  assign _04310_ = sel_oi_one_hot_i[163] & i[56];
  assign _04311_ = _04310_ | _04309_;
  assign _04312_ = _04311_ | _04308_;
  assign _04313_ = sel_oi_one_hot_i[164] & i[72];
  assign _04314_ = sel_oi_one_hot_i[165] & i[88];
  assign _04315_ = _04314_ | _04313_;
  assign _04316_ = sel_oi_one_hot_i[166] & i[104];
  assign _04317_ = sel_oi_one_hot_i[167] & i[120];
  assign _04318_ = _04317_ | _04316_;
  assign _04319_ = _04318_ | _04315_;
  assign _04320_ = _04319_ | _04312_;
  assign _04321_ = sel_oi_one_hot_i[168] & i[136];
  assign _04322_ = sel_oi_one_hot_i[169] & i[152];
  assign _04323_ = _04322_ | _04321_;
  assign _04324_ = sel_oi_one_hot_i[170] & i[168];
  assign _04325_ = sel_oi_one_hot_i[171] & i[184];
  assign _04326_ = _04325_ | _04324_;
  assign _04327_ = _04326_ | _04323_;
  assign _04328_ = sel_oi_one_hot_i[172] & i[200];
  assign _04329_ = sel_oi_one_hot_i[173] & i[216];
  assign _04330_ = _04329_ | _04328_;
  assign _04331_ = sel_oi_one_hot_i[174] & i[232];
  assign _04332_ = sel_oi_one_hot_i[175] & i[248];
  assign _04333_ = _04332_ | _04331_;
  assign _04334_ = _04333_ | _04330_;
  assign _04335_ = _04334_ | _04327_;
  assign o[168] = _04335_ | _04320_;
  assign _04336_ = sel_oi_one_hot_i[160] & i[7];
  assign _04337_ = sel_oi_one_hot_i[161] & i[23];
  assign _04338_ = _04337_ | _04336_;
  assign _04339_ = sel_oi_one_hot_i[162] & i[39];
  assign _04340_ = sel_oi_one_hot_i[163] & i[55];
  assign _04341_ = _04340_ | _04339_;
  assign _04342_ = _04341_ | _04338_;
  assign _04343_ = sel_oi_one_hot_i[164] & i[71];
  assign _04344_ = sel_oi_one_hot_i[165] & i[87];
  assign _04345_ = _04344_ | _04343_;
  assign _04346_ = sel_oi_one_hot_i[166] & i[103];
  assign _04347_ = sel_oi_one_hot_i[167] & i[119];
  assign _04348_ = _04347_ | _04346_;
  assign _04349_ = _04348_ | _04345_;
  assign _04350_ = _04349_ | _04342_;
  assign _04351_ = sel_oi_one_hot_i[168] & i[135];
  assign _04352_ = sel_oi_one_hot_i[169] & i[151];
  assign _04353_ = _04352_ | _04351_;
  assign _04354_ = sel_oi_one_hot_i[170] & i[167];
  assign _04355_ = sel_oi_one_hot_i[171] & i[183];
  assign _04356_ = _04355_ | _04354_;
  assign _04357_ = _04356_ | _04353_;
  assign _04358_ = sel_oi_one_hot_i[172] & i[199];
  assign _04359_ = sel_oi_one_hot_i[173] & i[215];
  assign _04360_ = _04359_ | _04358_;
  assign _04361_ = sel_oi_one_hot_i[174] & i[231];
  assign _04362_ = sel_oi_one_hot_i[175] & i[247];
  assign _04363_ = _04362_ | _04361_;
  assign _04364_ = _04363_ | _04360_;
  assign _04365_ = _04364_ | _04357_;
  assign o[167] = _04365_ | _04350_;
  assign _04366_ = sel_oi_one_hot_i[160] & i[6];
  assign _04367_ = sel_oi_one_hot_i[161] & i[22];
  assign _04368_ = _04367_ | _04366_;
  assign _04369_ = sel_oi_one_hot_i[162] & i[38];
  assign _04370_ = sel_oi_one_hot_i[163] & i[54];
  assign _04371_ = _04370_ | _04369_;
  assign _04372_ = _04371_ | _04368_;
  assign _04373_ = sel_oi_one_hot_i[164] & i[70];
  assign _04374_ = sel_oi_one_hot_i[165] & i[86];
  assign _04375_ = _04374_ | _04373_;
  assign _04376_ = sel_oi_one_hot_i[166] & i[102];
  assign _04377_ = sel_oi_one_hot_i[167] & i[118];
  assign _04378_ = _04377_ | _04376_;
  assign _04379_ = _04378_ | _04375_;
  assign _04380_ = _04379_ | _04372_;
  assign _04381_ = sel_oi_one_hot_i[168] & i[134];
  assign _04382_ = sel_oi_one_hot_i[169] & i[150];
  assign _04383_ = _04382_ | _04381_;
  assign _04384_ = sel_oi_one_hot_i[170] & i[166];
  assign _04385_ = sel_oi_one_hot_i[171] & i[182];
  assign _04386_ = _04385_ | _04384_;
  assign _04387_ = _04386_ | _04383_;
  assign _04388_ = sel_oi_one_hot_i[172] & i[198];
  assign _04389_ = sel_oi_one_hot_i[173] & i[214];
  assign _04390_ = _04389_ | _04388_;
  assign _04391_ = sel_oi_one_hot_i[174] & i[230];
  assign _04392_ = sel_oi_one_hot_i[175] & i[246];
  assign _04393_ = _04392_ | _04391_;
  assign _04394_ = _04393_ | _04390_;
  assign _04395_ = _04394_ | _04387_;
  assign o[166] = _04395_ | _04380_;
  assign _04396_ = sel_oi_one_hot_i[160] & i[5];
  assign _04397_ = sel_oi_one_hot_i[161] & i[21];
  assign _04398_ = _04397_ | _04396_;
  assign _04399_ = sel_oi_one_hot_i[162] & i[37];
  assign _04400_ = sel_oi_one_hot_i[163] & i[53];
  assign _04401_ = _04400_ | _04399_;
  assign _04402_ = _04401_ | _04398_;
  assign _04403_ = sel_oi_one_hot_i[164] & i[69];
  assign _04404_ = sel_oi_one_hot_i[165] & i[85];
  assign _04405_ = _04404_ | _04403_;
  assign _04406_ = sel_oi_one_hot_i[166] & i[101];
  assign _04407_ = sel_oi_one_hot_i[167] & i[117];
  assign _04408_ = _04407_ | _04406_;
  assign _04409_ = _04408_ | _04405_;
  assign _04410_ = _04409_ | _04402_;
  assign _04411_ = sel_oi_one_hot_i[168] & i[133];
  assign _04412_ = sel_oi_one_hot_i[169] & i[149];
  assign _04413_ = _04412_ | _04411_;
  assign _04414_ = sel_oi_one_hot_i[170] & i[165];
  assign _04415_ = sel_oi_one_hot_i[171] & i[181];
  assign _04416_ = _04415_ | _04414_;
  assign _04417_ = _04416_ | _04413_;
  assign _04418_ = sel_oi_one_hot_i[172] & i[197];
  assign _04419_ = sel_oi_one_hot_i[173] & i[213];
  assign _04420_ = _04419_ | _04418_;
  assign _04421_ = sel_oi_one_hot_i[174] & i[229];
  assign _04422_ = sel_oi_one_hot_i[175] & i[245];
  assign _04423_ = _04422_ | _04421_;
  assign _04424_ = _04423_ | _04420_;
  assign _04425_ = _04424_ | _04417_;
  assign o[165] = _04425_ | _04410_;
  assign _04426_ = sel_oi_one_hot_i[160] & i[4];
  assign _04427_ = sel_oi_one_hot_i[161] & i[20];
  assign _04428_ = _04427_ | _04426_;
  assign _04429_ = sel_oi_one_hot_i[162] & i[36];
  assign _04430_ = sel_oi_one_hot_i[163] & i[52];
  assign _04431_ = _04430_ | _04429_;
  assign _04432_ = _04431_ | _04428_;
  assign _04433_ = sel_oi_one_hot_i[164] & i[68];
  assign _04434_ = sel_oi_one_hot_i[165] & i[84];
  assign _04435_ = _04434_ | _04433_;
  assign _04436_ = sel_oi_one_hot_i[166] & i[100];
  assign _04437_ = sel_oi_one_hot_i[167] & i[116];
  assign _04438_ = _04437_ | _04436_;
  assign _04439_ = _04438_ | _04435_;
  assign _04440_ = _04439_ | _04432_;
  assign _04441_ = sel_oi_one_hot_i[168] & i[132];
  assign _04442_ = sel_oi_one_hot_i[169] & i[148];
  assign _04443_ = _04442_ | _04441_;
  assign _04444_ = sel_oi_one_hot_i[170] & i[164];
  assign _04445_ = sel_oi_one_hot_i[171] & i[180];
  assign _04446_ = _04445_ | _04444_;
  assign _04447_ = _04446_ | _04443_;
  assign _04448_ = sel_oi_one_hot_i[172] & i[196];
  assign _04449_ = sel_oi_one_hot_i[173] & i[212];
  assign _04450_ = _04449_ | _04448_;
  assign _04451_ = sel_oi_one_hot_i[174] & i[228];
  assign _04452_ = sel_oi_one_hot_i[175] & i[244];
  assign _04453_ = _04452_ | _04451_;
  assign _04454_ = _04453_ | _04450_;
  assign _04455_ = _04454_ | _04447_;
  assign o[164] = _04455_ | _04440_;
  assign _04456_ = sel_oi_one_hot_i[160] & i[3];
  assign _04457_ = sel_oi_one_hot_i[161] & i[19];
  assign _04458_ = _04457_ | _04456_;
  assign _04459_ = sel_oi_one_hot_i[162] & i[35];
  assign _04460_ = sel_oi_one_hot_i[163] & i[51];
  assign _04461_ = _04460_ | _04459_;
  assign _04462_ = _04461_ | _04458_;
  assign _04463_ = sel_oi_one_hot_i[164] & i[67];
  assign _04464_ = sel_oi_one_hot_i[165] & i[83];
  assign _04465_ = _04464_ | _04463_;
  assign _04466_ = sel_oi_one_hot_i[166] & i[99];
  assign _04467_ = sel_oi_one_hot_i[167] & i[115];
  assign _04468_ = _04467_ | _04466_;
  assign _04469_ = _04468_ | _04465_;
  assign _04470_ = _04469_ | _04462_;
  assign _04471_ = sel_oi_one_hot_i[168] & i[131];
  assign _04472_ = sel_oi_one_hot_i[169] & i[147];
  assign _04473_ = _04472_ | _04471_;
  assign _04474_ = sel_oi_one_hot_i[170] & i[163];
  assign _04475_ = sel_oi_one_hot_i[171] & i[179];
  assign _04476_ = _04475_ | _04474_;
  assign _04477_ = _04476_ | _04473_;
  assign _04478_ = sel_oi_one_hot_i[172] & i[195];
  assign _04479_ = sel_oi_one_hot_i[173] & i[211];
  assign _04480_ = _04479_ | _04478_;
  assign _04481_ = sel_oi_one_hot_i[174] & i[227];
  assign _04482_ = sel_oi_one_hot_i[175] & i[243];
  assign _04483_ = _04482_ | _04481_;
  assign _04484_ = _04483_ | _04480_;
  assign _04485_ = _04484_ | _04477_;
  assign o[163] = _04485_ | _04470_;
  assign _04486_ = sel_oi_one_hot_i[160] & i[2];
  assign _04487_ = sel_oi_one_hot_i[161] & i[18];
  assign _04488_ = _04487_ | _04486_;
  assign _04489_ = sel_oi_one_hot_i[162] & i[34];
  assign _04490_ = sel_oi_one_hot_i[163] & i[50];
  assign _04491_ = _04490_ | _04489_;
  assign _04492_ = _04491_ | _04488_;
  assign _04493_ = sel_oi_one_hot_i[164] & i[66];
  assign _04494_ = sel_oi_one_hot_i[165] & i[82];
  assign _04495_ = _04494_ | _04493_;
  assign _04496_ = sel_oi_one_hot_i[166] & i[98];
  assign _04497_ = sel_oi_one_hot_i[167] & i[114];
  assign _04498_ = _04497_ | _04496_;
  assign _04499_ = _04498_ | _04495_;
  assign _04500_ = _04499_ | _04492_;
  assign _04501_ = sel_oi_one_hot_i[168] & i[130];
  assign _04502_ = sel_oi_one_hot_i[169] & i[146];
  assign _04503_ = _04502_ | _04501_;
  assign _04504_ = sel_oi_one_hot_i[170] & i[162];
  assign _04505_ = sel_oi_one_hot_i[171] & i[178];
  assign _04506_ = _04505_ | _04504_;
  assign _04507_ = _04506_ | _04503_;
  assign _04508_ = sel_oi_one_hot_i[172] & i[194];
  assign _04509_ = sel_oi_one_hot_i[173] & i[210];
  assign _04510_ = _04509_ | _04508_;
  assign _04511_ = sel_oi_one_hot_i[174] & i[226];
  assign _04512_ = sel_oi_one_hot_i[175] & i[242];
  assign _04513_ = _04512_ | _04511_;
  assign _04514_ = _04513_ | _04510_;
  assign _04515_ = _04514_ | _04507_;
  assign o[162] = _04515_ | _04500_;
  assign _04516_ = sel_oi_one_hot_i[160] & i[1];
  assign _04517_ = sel_oi_one_hot_i[161] & i[17];
  assign _04518_ = _04517_ | _04516_;
  assign _04519_ = sel_oi_one_hot_i[162] & i[33];
  assign _04520_ = sel_oi_one_hot_i[163] & i[49];
  assign _04521_ = _04520_ | _04519_;
  assign _04522_ = _04521_ | _04518_;
  assign _04523_ = sel_oi_one_hot_i[164] & i[65];
  assign _04524_ = sel_oi_one_hot_i[165] & i[81];
  assign _04525_ = _04524_ | _04523_;
  assign _04526_ = sel_oi_one_hot_i[166] & i[97];
  assign _04527_ = sel_oi_one_hot_i[167] & i[113];
  assign _04528_ = _04527_ | _04526_;
  assign _04529_ = _04528_ | _04525_;
  assign _04530_ = _04529_ | _04522_;
  assign _04531_ = sel_oi_one_hot_i[168] & i[129];
  assign _04532_ = sel_oi_one_hot_i[169] & i[145];
  assign _04533_ = _04532_ | _04531_;
  assign _04534_ = sel_oi_one_hot_i[170] & i[161];
  assign _04535_ = sel_oi_one_hot_i[171] & i[177];
  assign _04536_ = _04535_ | _04534_;
  assign _04537_ = _04536_ | _04533_;
  assign _04538_ = sel_oi_one_hot_i[172] & i[193];
  assign _04539_ = sel_oi_one_hot_i[173] & i[209];
  assign _04540_ = _04539_ | _04538_;
  assign _04541_ = sel_oi_one_hot_i[174] & i[225];
  assign _04542_ = sel_oi_one_hot_i[175] & i[241];
  assign _04543_ = _04542_ | _04541_;
  assign _04544_ = _04543_ | _04540_;
  assign _04545_ = _04544_ | _04537_;
  assign o[161] = _04545_ | _04530_;
  assign _04546_ = sel_oi_one_hot_i[160] & i[0];
  assign _04547_ = sel_oi_one_hot_i[161] & i[16];
  assign _04548_ = _04547_ | _04546_;
  assign _04549_ = sel_oi_one_hot_i[162] & i[32];
  assign _04550_ = sel_oi_one_hot_i[163] & i[48];
  assign _04551_ = _04550_ | _04549_;
  assign _04552_ = _04551_ | _04548_;
  assign _04553_ = sel_oi_one_hot_i[164] & i[64];
  assign _04554_ = sel_oi_one_hot_i[165] & i[80];
  assign _04555_ = _04554_ | _04553_;
  assign _04556_ = sel_oi_one_hot_i[166] & i[96];
  assign _04557_ = sel_oi_one_hot_i[167] & i[112];
  assign _04558_ = _04557_ | _04556_;
  assign _04559_ = _04558_ | _04555_;
  assign _04560_ = _04559_ | _04552_;
  assign _04561_ = sel_oi_one_hot_i[168] & i[128];
  assign _04562_ = sel_oi_one_hot_i[169] & i[144];
  assign _04563_ = _04562_ | _04561_;
  assign _04564_ = sel_oi_one_hot_i[170] & i[160];
  assign _04565_ = sel_oi_one_hot_i[171] & i[176];
  assign _04566_ = _04565_ | _04564_;
  assign _04567_ = _04566_ | _04563_;
  assign _04568_ = sel_oi_one_hot_i[172] & i[192];
  assign _04569_ = sel_oi_one_hot_i[173] & i[208];
  assign _04570_ = _04569_ | _04568_;
  assign _04571_ = sel_oi_one_hot_i[174] & i[224];
  assign _04572_ = sel_oi_one_hot_i[175] & i[240];
  assign _04573_ = _04572_ | _04571_;
  assign _04574_ = _04573_ | _04570_;
  assign _04575_ = _04574_ | _04567_;
  assign o[160] = _04575_ | _04560_;
  assign _04576_ = sel_oi_one_hot_i[176] & i[15];
  assign _04577_ = sel_oi_one_hot_i[177] & i[31];
  assign _04578_ = _04577_ | _04576_;
  assign _04579_ = sel_oi_one_hot_i[178] & i[47];
  assign _04580_ = sel_oi_one_hot_i[179] & i[63];
  assign _04581_ = _04580_ | _04579_;
  assign _04582_ = _04581_ | _04578_;
  assign _04583_ = sel_oi_one_hot_i[180] & i[79];
  assign _04584_ = sel_oi_one_hot_i[181] & i[95];
  assign _04585_ = _04584_ | _04583_;
  assign _04586_ = sel_oi_one_hot_i[182] & i[111];
  assign _04587_ = sel_oi_one_hot_i[183] & i[127];
  assign _04588_ = _04587_ | _04586_;
  assign _04589_ = _04588_ | _04585_;
  assign _04590_ = _04589_ | _04582_;
  assign _04591_ = sel_oi_one_hot_i[184] & i[143];
  assign _04592_ = sel_oi_one_hot_i[185] & i[159];
  assign _04593_ = _04592_ | _04591_;
  assign _04594_ = sel_oi_one_hot_i[186] & i[175];
  assign _04595_ = sel_oi_one_hot_i[187] & i[191];
  assign _04596_ = _04595_ | _04594_;
  assign _04597_ = _04596_ | _04593_;
  assign _04598_ = sel_oi_one_hot_i[188] & i[207];
  assign _04599_ = sel_oi_one_hot_i[189] & i[223];
  assign _04600_ = _04599_ | _04598_;
  assign _04601_ = sel_oi_one_hot_i[190] & i[239];
  assign _04602_ = sel_oi_one_hot_i[191] & i[255];
  assign _04603_ = _04602_ | _04601_;
  assign _04604_ = _04603_ | _04600_;
  assign _04605_ = _04604_ | _04597_;
  assign o[191] = _04605_ | _04590_;
  assign _04606_ = sel_oi_one_hot_i[176] & i[14];
  assign _04607_ = sel_oi_one_hot_i[177] & i[30];
  assign _04608_ = _04607_ | _04606_;
  assign _04609_ = sel_oi_one_hot_i[178] & i[46];
  assign _04610_ = sel_oi_one_hot_i[179] & i[62];
  assign _04611_ = _04610_ | _04609_;
  assign _04612_ = _04611_ | _04608_;
  assign _04613_ = sel_oi_one_hot_i[180] & i[78];
  assign _04614_ = sel_oi_one_hot_i[181] & i[94];
  assign _04615_ = _04614_ | _04613_;
  assign _04616_ = sel_oi_one_hot_i[182] & i[110];
  assign _04617_ = sel_oi_one_hot_i[183] & i[126];
  assign _04618_ = _04617_ | _04616_;
  assign _04619_ = _04618_ | _04615_;
  assign _04620_ = _04619_ | _04612_;
  assign _04621_ = sel_oi_one_hot_i[184] & i[142];
  assign _04622_ = sel_oi_one_hot_i[185] & i[158];
  assign _04623_ = _04622_ | _04621_;
  assign _04624_ = sel_oi_one_hot_i[186] & i[174];
  assign _04625_ = sel_oi_one_hot_i[187] & i[190];
  assign _04626_ = _04625_ | _04624_;
  assign _04627_ = _04626_ | _04623_;
  assign _04628_ = sel_oi_one_hot_i[188] & i[206];
  assign _04629_ = sel_oi_one_hot_i[189] & i[222];
  assign _04630_ = _04629_ | _04628_;
  assign _04631_ = sel_oi_one_hot_i[190] & i[238];
  assign _04632_ = sel_oi_one_hot_i[191] & i[254];
  assign _04633_ = _04632_ | _04631_;
  assign _04634_ = _04633_ | _04630_;
  assign _04635_ = _04634_ | _04627_;
  assign o[190] = _04635_ | _04620_;
  assign _04636_ = sel_oi_one_hot_i[176] & i[13];
  assign _04637_ = sel_oi_one_hot_i[177] & i[29];
  assign _04638_ = _04637_ | _04636_;
  assign _04639_ = sel_oi_one_hot_i[178] & i[45];
  assign _04640_ = sel_oi_one_hot_i[179] & i[61];
  assign _04641_ = _04640_ | _04639_;
  assign _04642_ = _04641_ | _04638_;
  assign _04643_ = sel_oi_one_hot_i[180] & i[77];
  assign _04644_ = sel_oi_one_hot_i[181] & i[93];
  assign _04645_ = _04644_ | _04643_;
  assign _04646_ = sel_oi_one_hot_i[182] & i[109];
  assign _04647_ = sel_oi_one_hot_i[183] & i[125];
  assign _04648_ = _04647_ | _04646_;
  assign _04649_ = _04648_ | _04645_;
  assign _04650_ = _04649_ | _04642_;
  assign _04651_ = sel_oi_one_hot_i[184] & i[141];
  assign _04652_ = sel_oi_one_hot_i[185] & i[157];
  assign _04653_ = _04652_ | _04651_;
  assign _04654_ = sel_oi_one_hot_i[186] & i[173];
  assign _04655_ = sel_oi_one_hot_i[187] & i[189];
  assign _04656_ = _04655_ | _04654_;
  assign _04657_ = _04656_ | _04653_;
  assign _04658_ = sel_oi_one_hot_i[188] & i[205];
  assign _04659_ = sel_oi_one_hot_i[189] & i[221];
  assign _04660_ = _04659_ | _04658_;
  assign _04661_ = sel_oi_one_hot_i[190] & i[237];
  assign _04662_ = sel_oi_one_hot_i[191] & i[253];
  assign _04663_ = _04662_ | _04661_;
  assign _04664_ = _04663_ | _04660_;
  assign _04665_ = _04664_ | _04657_;
  assign o[189] = _04665_ | _04650_;
  assign _04666_ = sel_oi_one_hot_i[176] & i[12];
  assign _04667_ = sel_oi_one_hot_i[177] & i[28];
  assign _04668_ = _04667_ | _04666_;
  assign _04669_ = sel_oi_one_hot_i[178] & i[44];
  assign _04670_ = sel_oi_one_hot_i[179] & i[60];
  assign _04671_ = _04670_ | _04669_;
  assign _04672_ = _04671_ | _04668_;
  assign _04673_ = sel_oi_one_hot_i[180] & i[76];
  assign _04674_ = sel_oi_one_hot_i[181] & i[92];
  assign _04675_ = _04674_ | _04673_;
  assign _04676_ = sel_oi_one_hot_i[182] & i[108];
  assign _04677_ = sel_oi_one_hot_i[183] & i[124];
  assign _04678_ = _04677_ | _04676_;
  assign _04679_ = _04678_ | _04675_;
  assign _04680_ = _04679_ | _04672_;
  assign _04681_ = sel_oi_one_hot_i[184] & i[140];
  assign _04682_ = sel_oi_one_hot_i[185] & i[156];
  assign _04683_ = _04682_ | _04681_;
  assign _04684_ = sel_oi_one_hot_i[186] & i[172];
  assign _04685_ = sel_oi_one_hot_i[187] & i[188];
  assign _04686_ = _04685_ | _04684_;
  assign _04687_ = _04686_ | _04683_;
  assign _04688_ = sel_oi_one_hot_i[188] & i[204];
  assign _04689_ = sel_oi_one_hot_i[189] & i[220];
  assign _04690_ = _04689_ | _04688_;
  assign _04691_ = sel_oi_one_hot_i[190] & i[236];
  assign _04692_ = sel_oi_one_hot_i[191] & i[252];
  assign _04693_ = _04692_ | _04691_;
  assign _04694_ = _04693_ | _04690_;
  assign _04695_ = _04694_ | _04687_;
  assign o[188] = _04695_ | _04680_;
  assign _04696_ = sel_oi_one_hot_i[176] & i[11];
  assign _04697_ = sel_oi_one_hot_i[177] & i[27];
  assign _04698_ = _04697_ | _04696_;
  assign _04699_ = sel_oi_one_hot_i[178] & i[43];
  assign _04700_ = sel_oi_one_hot_i[179] & i[59];
  assign _04701_ = _04700_ | _04699_;
  assign _04702_ = _04701_ | _04698_;
  assign _04703_ = sel_oi_one_hot_i[180] & i[75];
  assign _04704_ = sel_oi_one_hot_i[181] & i[91];
  assign _04705_ = _04704_ | _04703_;
  assign _04706_ = sel_oi_one_hot_i[182] & i[107];
  assign _04707_ = sel_oi_one_hot_i[183] & i[123];
  assign _04708_ = _04707_ | _04706_;
  assign _04709_ = _04708_ | _04705_;
  assign _04710_ = _04709_ | _04702_;
  assign _04711_ = sel_oi_one_hot_i[184] & i[139];
  assign _04712_ = sel_oi_one_hot_i[185] & i[155];
  assign _04713_ = _04712_ | _04711_;
  assign _04714_ = sel_oi_one_hot_i[186] & i[171];
  assign _04715_ = sel_oi_one_hot_i[187] & i[187];
  assign _04716_ = _04715_ | _04714_;
  assign _04717_ = _04716_ | _04713_;
  assign _04718_ = sel_oi_one_hot_i[188] & i[203];
  assign _04719_ = sel_oi_one_hot_i[189] & i[219];
  assign _04720_ = _04719_ | _04718_;
  assign _04721_ = sel_oi_one_hot_i[190] & i[235];
  assign _04722_ = sel_oi_one_hot_i[191] & i[251];
  assign _04723_ = _04722_ | _04721_;
  assign _04724_ = _04723_ | _04720_;
  assign _04725_ = _04724_ | _04717_;
  assign o[187] = _04725_ | _04710_;
  assign _04726_ = sel_oi_one_hot_i[176] & i[10];
  assign _04727_ = sel_oi_one_hot_i[177] & i[26];
  assign _04728_ = _04727_ | _04726_;
  assign _04729_ = sel_oi_one_hot_i[178] & i[42];
  assign _04730_ = sel_oi_one_hot_i[179] & i[58];
  assign _04731_ = _04730_ | _04729_;
  assign _04732_ = _04731_ | _04728_;
  assign _04733_ = sel_oi_one_hot_i[180] & i[74];
  assign _04734_ = sel_oi_one_hot_i[181] & i[90];
  assign _04735_ = _04734_ | _04733_;
  assign _04736_ = sel_oi_one_hot_i[182] & i[106];
  assign _04737_ = sel_oi_one_hot_i[183] & i[122];
  assign _04738_ = _04737_ | _04736_;
  assign _04739_ = _04738_ | _04735_;
  assign _04740_ = _04739_ | _04732_;
  assign _04741_ = sel_oi_one_hot_i[184] & i[138];
  assign _04742_ = sel_oi_one_hot_i[185] & i[154];
  assign _04743_ = _04742_ | _04741_;
  assign _04744_ = sel_oi_one_hot_i[186] & i[170];
  assign _04745_ = sel_oi_one_hot_i[187] & i[186];
  assign _04746_ = _04745_ | _04744_;
  assign _04747_ = _04746_ | _04743_;
  assign _04748_ = sel_oi_one_hot_i[188] & i[202];
  assign _04749_ = sel_oi_one_hot_i[189] & i[218];
  assign _04750_ = _04749_ | _04748_;
  assign _04751_ = sel_oi_one_hot_i[190] & i[234];
  assign _04752_ = sel_oi_one_hot_i[191] & i[250];
  assign _04753_ = _04752_ | _04751_;
  assign _04754_ = _04753_ | _04750_;
  assign _04755_ = _04754_ | _04747_;
  assign o[186] = _04755_ | _04740_;
  assign _04756_ = sel_oi_one_hot_i[176] & i[9];
  assign _04757_ = sel_oi_one_hot_i[177] & i[25];
  assign _04758_ = _04757_ | _04756_;
  assign _04759_ = sel_oi_one_hot_i[178] & i[41];
  assign _04760_ = sel_oi_one_hot_i[179] & i[57];
  assign _04761_ = _04760_ | _04759_;
  assign _04762_ = _04761_ | _04758_;
  assign _04763_ = sel_oi_one_hot_i[180] & i[73];
  assign _04764_ = sel_oi_one_hot_i[181] & i[89];
  assign _04765_ = _04764_ | _04763_;
  assign _04766_ = sel_oi_one_hot_i[182] & i[105];
  assign _04767_ = sel_oi_one_hot_i[183] & i[121];
  assign _04768_ = _04767_ | _04766_;
  assign _04769_ = _04768_ | _04765_;
  assign _04770_ = _04769_ | _04762_;
  assign _04771_ = sel_oi_one_hot_i[184] & i[137];
  assign _04772_ = sel_oi_one_hot_i[185] & i[153];
  assign _04773_ = _04772_ | _04771_;
  assign _04774_ = sel_oi_one_hot_i[186] & i[169];
  assign _04775_ = sel_oi_one_hot_i[187] & i[185];
  assign _04776_ = _04775_ | _04774_;
  assign _04777_ = _04776_ | _04773_;
  assign _04778_ = sel_oi_one_hot_i[188] & i[201];
  assign _04779_ = sel_oi_one_hot_i[189] & i[217];
  assign _04780_ = _04779_ | _04778_;
  assign _04781_ = sel_oi_one_hot_i[190] & i[233];
  assign _04782_ = sel_oi_one_hot_i[191] & i[249];
  assign _04783_ = _04782_ | _04781_;
  assign _04784_ = _04783_ | _04780_;
  assign _04785_ = _04784_ | _04777_;
  assign o[185] = _04785_ | _04770_;
  assign _04786_ = sel_oi_one_hot_i[176] & i[8];
  assign _04787_ = sel_oi_one_hot_i[177] & i[24];
  assign _04788_ = _04787_ | _04786_;
  assign _04789_ = sel_oi_one_hot_i[178] & i[40];
  assign _04790_ = sel_oi_one_hot_i[179] & i[56];
  assign _04791_ = _04790_ | _04789_;
  assign _04792_ = _04791_ | _04788_;
  assign _04793_ = sel_oi_one_hot_i[180] & i[72];
  assign _04794_ = sel_oi_one_hot_i[181] & i[88];
  assign _04795_ = _04794_ | _04793_;
  assign _04796_ = sel_oi_one_hot_i[182] & i[104];
  assign _04797_ = sel_oi_one_hot_i[183] & i[120];
  assign _04798_ = _04797_ | _04796_;
  assign _04799_ = _04798_ | _04795_;
  assign _04800_ = _04799_ | _04792_;
  assign _04801_ = sel_oi_one_hot_i[184] & i[136];
  assign _04802_ = sel_oi_one_hot_i[185] & i[152];
  assign _04803_ = _04802_ | _04801_;
  assign _04804_ = sel_oi_one_hot_i[186] & i[168];
  assign _04805_ = sel_oi_one_hot_i[187] & i[184];
  assign _04806_ = _04805_ | _04804_;
  assign _04807_ = _04806_ | _04803_;
  assign _04808_ = sel_oi_one_hot_i[188] & i[200];
  assign _04809_ = sel_oi_one_hot_i[189] & i[216];
  assign _04810_ = _04809_ | _04808_;
  assign _04811_ = sel_oi_one_hot_i[190] & i[232];
  assign _04812_ = sel_oi_one_hot_i[191] & i[248];
  assign _04813_ = _04812_ | _04811_;
  assign _04814_ = _04813_ | _04810_;
  assign _04815_ = _04814_ | _04807_;
  assign o[184] = _04815_ | _04800_;
  assign _04816_ = sel_oi_one_hot_i[176] & i[7];
  assign _04817_ = sel_oi_one_hot_i[177] & i[23];
  assign _04818_ = _04817_ | _04816_;
  assign _04819_ = sel_oi_one_hot_i[178] & i[39];
  assign _04820_ = sel_oi_one_hot_i[179] & i[55];
  assign _04821_ = _04820_ | _04819_;
  assign _04822_ = _04821_ | _04818_;
  assign _04823_ = sel_oi_one_hot_i[180] & i[71];
  assign _04824_ = sel_oi_one_hot_i[181] & i[87];
  assign _04825_ = _04824_ | _04823_;
  assign _04826_ = sel_oi_one_hot_i[182] & i[103];
  assign _04827_ = sel_oi_one_hot_i[183] & i[119];
  assign _04828_ = _04827_ | _04826_;
  assign _04829_ = _04828_ | _04825_;
  assign _04830_ = _04829_ | _04822_;
  assign _04831_ = sel_oi_one_hot_i[184] & i[135];
  assign _04832_ = sel_oi_one_hot_i[185] & i[151];
  assign _04833_ = _04832_ | _04831_;
  assign _04834_ = sel_oi_one_hot_i[186] & i[167];
  assign _04835_ = sel_oi_one_hot_i[187] & i[183];
  assign _04836_ = _04835_ | _04834_;
  assign _04837_ = _04836_ | _04833_;
  assign _04838_ = sel_oi_one_hot_i[188] & i[199];
  assign _04839_ = sel_oi_one_hot_i[189] & i[215];
  assign _04840_ = _04839_ | _04838_;
  assign _04841_ = sel_oi_one_hot_i[190] & i[231];
  assign _04842_ = sel_oi_one_hot_i[191] & i[247];
  assign _04843_ = _04842_ | _04841_;
  assign _04844_ = _04843_ | _04840_;
  assign _04845_ = _04844_ | _04837_;
  assign o[183] = _04845_ | _04830_;
  assign _04846_ = sel_oi_one_hot_i[176] & i[6];
  assign _04847_ = sel_oi_one_hot_i[177] & i[22];
  assign _04848_ = _04847_ | _04846_;
  assign _04849_ = sel_oi_one_hot_i[178] & i[38];
  assign _04850_ = sel_oi_one_hot_i[179] & i[54];
  assign _04851_ = _04850_ | _04849_;
  assign _04852_ = _04851_ | _04848_;
  assign _04853_ = sel_oi_one_hot_i[180] & i[70];
  assign _04854_ = sel_oi_one_hot_i[181] & i[86];
  assign _04855_ = _04854_ | _04853_;
  assign _04856_ = sel_oi_one_hot_i[182] & i[102];
  assign _04857_ = sel_oi_one_hot_i[183] & i[118];
  assign _04858_ = _04857_ | _04856_;
  assign _04859_ = _04858_ | _04855_;
  assign _04860_ = _04859_ | _04852_;
  assign _04861_ = sel_oi_one_hot_i[184] & i[134];
  assign _04862_ = sel_oi_one_hot_i[185] & i[150];
  assign _04863_ = _04862_ | _04861_;
  assign _04864_ = sel_oi_one_hot_i[186] & i[166];
  assign _04865_ = sel_oi_one_hot_i[187] & i[182];
  assign _04866_ = _04865_ | _04864_;
  assign _04867_ = _04866_ | _04863_;
  assign _04868_ = sel_oi_one_hot_i[188] & i[198];
  assign _04869_ = sel_oi_one_hot_i[189] & i[214];
  assign _04870_ = _04869_ | _04868_;
  assign _04871_ = sel_oi_one_hot_i[190] & i[230];
  assign _04872_ = sel_oi_one_hot_i[191] & i[246];
  assign _04873_ = _04872_ | _04871_;
  assign _04874_ = _04873_ | _04870_;
  assign _04875_ = _04874_ | _04867_;
  assign o[182] = _04875_ | _04860_;
  assign _04876_ = sel_oi_one_hot_i[176] & i[5];
  assign _04877_ = sel_oi_one_hot_i[177] & i[21];
  assign _04878_ = _04877_ | _04876_;
  assign _04879_ = sel_oi_one_hot_i[178] & i[37];
  assign _04880_ = sel_oi_one_hot_i[179] & i[53];
  assign _04881_ = _04880_ | _04879_;
  assign _04882_ = _04881_ | _04878_;
  assign _04883_ = sel_oi_one_hot_i[180] & i[69];
  assign _04884_ = sel_oi_one_hot_i[181] & i[85];
  assign _04885_ = _04884_ | _04883_;
  assign _04886_ = sel_oi_one_hot_i[182] & i[101];
  assign _04887_ = sel_oi_one_hot_i[183] & i[117];
  assign _04888_ = _04887_ | _04886_;
  assign _04889_ = _04888_ | _04885_;
  assign _04890_ = _04889_ | _04882_;
  assign _04891_ = sel_oi_one_hot_i[184] & i[133];
  assign _04892_ = sel_oi_one_hot_i[185] & i[149];
  assign _04893_ = _04892_ | _04891_;
  assign _04894_ = sel_oi_one_hot_i[186] & i[165];
  assign _04895_ = sel_oi_one_hot_i[187] & i[181];
  assign _04896_ = _04895_ | _04894_;
  assign _04897_ = _04896_ | _04893_;
  assign _04898_ = sel_oi_one_hot_i[188] & i[197];
  assign _04899_ = sel_oi_one_hot_i[189] & i[213];
  assign _04900_ = _04899_ | _04898_;
  assign _04901_ = sel_oi_one_hot_i[190] & i[229];
  assign _04902_ = sel_oi_one_hot_i[191] & i[245];
  assign _04903_ = _04902_ | _04901_;
  assign _04904_ = _04903_ | _04900_;
  assign _04905_ = _04904_ | _04897_;
  assign o[181] = _04905_ | _04890_;
  assign _04906_ = sel_oi_one_hot_i[176] & i[4];
  assign _04907_ = sel_oi_one_hot_i[177] & i[20];
  assign _04908_ = _04907_ | _04906_;
  assign _04909_ = sel_oi_one_hot_i[178] & i[36];
  assign _04910_ = sel_oi_one_hot_i[179] & i[52];
  assign _04911_ = _04910_ | _04909_;
  assign _04912_ = _04911_ | _04908_;
  assign _04913_ = sel_oi_one_hot_i[180] & i[68];
  assign _04914_ = sel_oi_one_hot_i[181] & i[84];
  assign _04915_ = _04914_ | _04913_;
  assign _04916_ = sel_oi_one_hot_i[182] & i[100];
  assign _04917_ = sel_oi_one_hot_i[183] & i[116];
  assign _04918_ = _04917_ | _04916_;
  assign _04919_ = _04918_ | _04915_;
  assign _04920_ = _04919_ | _04912_;
  assign _04921_ = sel_oi_one_hot_i[184] & i[132];
  assign _04922_ = sel_oi_one_hot_i[185] & i[148];
  assign _04923_ = _04922_ | _04921_;
  assign _04924_ = sel_oi_one_hot_i[186] & i[164];
  assign _04925_ = sel_oi_one_hot_i[187] & i[180];
  assign _04926_ = _04925_ | _04924_;
  assign _04927_ = _04926_ | _04923_;
  assign _04928_ = sel_oi_one_hot_i[188] & i[196];
  assign _04929_ = sel_oi_one_hot_i[189] & i[212];
  assign _04930_ = _04929_ | _04928_;
  assign _04931_ = sel_oi_one_hot_i[190] & i[228];
  assign _04932_ = sel_oi_one_hot_i[191] & i[244];
  assign _04933_ = _04932_ | _04931_;
  assign _04934_ = _04933_ | _04930_;
  assign _04935_ = _04934_ | _04927_;
  assign o[180] = _04935_ | _04920_;
  assign _04936_ = sel_oi_one_hot_i[176] & i[3];
  assign _04937_ = sel_oi_one_hot_i[177] & i[19];
  assign _04938_ = _04937_ | _04936_;
  assign _04939_ = sel_oi_one_hot_i[178] & i[35];
  assign _04940_ = sel_oi_one_hot_i[179] & i[51];
  assign _04941_ = _04940_ | _04939_;
  assign _04942_ = _04941_ | _04938_;
  assign _04943_ = sel_oi_one_hot_i[180] & i[67];
  assign _04944_ = sel_oi_one_hot_i[181] & i[83];
  assign _04945_ = _04944_ | _04943_;
  assign _04946_ = sel_oi_one_hot_i[182] & i[99];
  assign _04947_ = sel_oi_one_hot_i[183] & i[115];
  assign _04948_ = _04947_ | _04946_;
  assign _04949_ = _04948_ | _04945_;
  assign _04950_ = _04949_ | _04942_;
  assign _04951_ = sel_oi_one_hot_i[184] & i[131];
  assign _04952_ = sel_oi_one_hot_i[185] & i[147];
  assign _04953_ = _04952_ | _04951_;
  assign _04954_ = sel_oi_one_hot_i[186] & i[163];
  assign _04955_ = sel_oi_one_hot_i[187] & i[179];
  assign _04956_ = _04955_ | _04954_;
  assign _04957_ = _04956_ | _04953_;
  assign _04958_ = sel_oi_one_hot_i[188] & i[195];
  assign _04959_ = sel_oi_one_hot_i[189] & i[211];
  assign _04960_ = _04959_ | _04958_;
  assign _04961_ = sel_oi_one_hot_i[190] & i[227];
  assign _04962_ = sel_oi_one_hot_i[191] & i[243];
  assign _04963_ = _04962_ | _04961_;
  assign _04964_ = _04963_ | _04960_;
  assign _04965_ = _04964_ | _04957_;
  assign o[179] = _04965_ | _04950_;
  assign _04966_ = sel_oi_one_hot_i[176] & i[2];
  assign _04967_ = sel_oi_one_hot_i[177] & i[18];
  assign _04968_ = _04967_ | _04966_;
  assign _04969_ = sel_oi_one_hot_i[178] & i[34];
  assign _04970_ = sel_oi_one_hot_i[179] & i[50];
  assign _04971_ = _04970_ | _04969_;
  assign _04972_ = _04971_ | _04968_;
  assign _04973_ = sel_oi_one_hot_i[180] & i[66];
  assign _04974_ = sel_oi_one_hot_i[181] & i[82];
  assign _04975_ = _04974_ | _04973_;
  assign _04976_ = sel_oi_one_hot_i[182] & i[98];
  assign _04977_ = sel_oi_one_hot_i[183] & i[114];
  assign _04978_ = _04977_ | _04976_;
  assign _04979_ = _04978_ | _04975_;
  assign _04980_ = _04979_ | _04972_;
  assign _04981_ = sel_oi_one_hot_i[184] & i[130];
  assign _04982_ = sel_oi_one_hot_i[185] & i[146];
  assign _04983_ = _04982_ | _04981_;
  assign _04984_ = sel_oi_one_hot_i[186] & i[162];
  assign _04985_ = sel_oi_one_hot_i[187] & i[178];
  assign _04986_ = _04985_ | _04984_;
  assign _04987_ = _04986_ | _04983_;
  assign _04988_ = sel_oi_one_hot_i[188] & i[194];
  assign _04989_ = sel_oi_one_hot_i[189] & i[210];
  assign _04990_ = _04989_ | _04988_;
  assign _04991_ = sel_oi_one_hot_i[190] & i[226];
  assign _04992_ = sel_oi_one_hot_i[191] & i[242];
  assign _04993_ = _04992_ | _04991_;
  assign _04994_ = _04993_ | _04990_;
  assign _04995_ = _04994_ | _04987_;
  assign o[178] = _04995_ | _04980_;
  assign _04996_ = sel_oi_one_hot_i[176] & i[1];
  assign _04997_ = sel_oi_one_hot_i[177] & i[17];
  assign _04998_ = _04997_ | _04996_;
  assign _04999_ = sel_oi_one_hot_i[178] & i[33];
  assign _05000_ = sel_oi_one_hot_i[179] & i[49];
  assign _05001_ = _05000_ | _04999_;
  assign _05002_ = _05001_ | _04998_;
  assign _05003_ = sel_oi_one_hot_i[180] & i[65];
  assign _05004_ = sel_oi_one_hot_i[181] & i[81];
  assign _05005_ = _05004_ | _05003_;
  assign _05006_ = sel_oi_one_hot_i[182] & i[97];
  assign _05007_ = sel_oi_one_hot_i[183] & i[113];
  assign _05008_ = _05007_ | _05006_;
  assign _05009_ = _05008_ | _05005_;
  assign _05010_ = _05009_ | _05002_;
  assign _05011_ = sel_oi_one_hot_i[184] & i[129];
  assign _05012_ = sel_oi_one_hot_i[185] & i[145];
  assign _05013_ = _05012_ | _05011_;
  assign _05014_ = sel_oi_one_hot_i[186] & i[161];
  assign _05015_ = sel_oi_one_hot_i[187] & i[177];
  assign _05016_ = _05015_ | _05014_;
  assign _05017_ = _05016_ | _05013_;
  assign _05018_ = sel_oi_one_hot_i[188] & i[193];
  assign _05019_ = sel_oi_one_hot_i[189] & i[209];
  assign _05020_ = _05019_ | _05018_;
  assign _05021_ = sel_oi_one_hot_i[190] & i[225];
  assign _05022_ = sel_oi_one_hot_i[191] & i[241];
  assign _05023_ = _05022_ | _05021_;
  assign _05024_ = _05023_ | _05020_;
  assign _05025_ = _05024_ | _05017_;
  assign o[177] = _05025_ | _05010_;
  assign _05026_ = sel_oi_one_hot_i[176] & i[0];
  assign _05027_ = sel_oi_one_hot_i[177] & i[16];
  assign _05028_ = _05027_ | _05026_;
  assign _05029_ = sel_oi_one_hot_i[178] & i[32];
  assign _05030_ = sel_oi_one_hot_i[179] & i[48];
  assign _05031_ = _05030_ | _05029_;
  assign _05032_ = _05031_ | _05028_;
  assign _05033_ = sel_oi_one_hot_i[180] & i[64];
  assign _05034_ = sel_oi_one_hot_i[181] & i[80];
  assign _05035_ = _05034_ | _05033_;
  assign _05036_ = sel_oi_one_hot_i[182] & i[96];
  assign _05037_ = sel_oi_one_hot_i[183] & i[112];
  assign _05038_ = _05037_ | _05036_;
  assign _05039_ = _05038_ | _05035_;
  assign _05040_ = _05039_ | _05032_;
  assign _05041_ = sel_oi_one_hot_i[184] & i[128];
  assign _05042_ = sel_oi_one_hot_i[185] & i[144];
  assign _05043_ = _05042_ | _05041_;
  assign _05044_ = sel_oi_one_hot_i[186] & i[160];
  assign _05045_ = sel_oi_one_hot_i[187] & i[176];
  assign _05046_ = _05045_ | _05044_;
  assign _05047_ = _05046_ | _05043_;
  assign _05048_ = sel_oi_one_hot_i[188] & i[192];
  assign _05049_ = sel_oi_one_hot_i[189] & i[208];
  assign _05050_ = _05049_ | _05048_;
  assign _05051_ = sel_oi_one_hot_i[190] & i[224];
  assign _05052_ = sel_oi_one_hot_i[191] & i[240];
  assign _05053_ = _05052_ | _05051_;
  assign _05054_ = _05053_ | _05050_;
  assign _05055_ = _05054_ | _05047_;
  assign o[176] = _05055_ | _05040_;
  assign _05056_ = sel_oi_one_hot_i[192] & i[15];
  assign _05057_ = sel_oi_one_hot_i[193] & i[31];
  assign _05058_ = _05057_ | _05056_;
  assign _05059_ = sel_oi_one_hot_i[194] & i[47];
  assign _05060_ = sel_oi_one_hot_i[195] & i[63];
  assign _05061_ = _05060_ | _05059_;
  assign _05062_ = _05061_ | _05058_;
  assign _05063_ = sel_oi_one_hot_i[196] & i[79];
  assign _05064_ = sel_oi_one_hot_i[197] & i[95];
  assign _05065_ = _05064_ | _05063_;
  assign _05066_ = sel_oi_one_hot_i[198] & i[111];
  assign _05067_ = sel_oi_one_hot_i[199] & i[127];
  assign _05068_ = _05067_ | _05066_;
  assign _05069_ = _05068_ | _05065_;
  assign _05070_ = _05069_ | _05062_;
  assign _05071_ = sel_oi_one_hot_i[200] & i[143];
  assign _05072_ = sel_oi_one_hot_i[201] & i[159];
  assign _05073_ = _05072_ | _05071_;
  assign _05074_ = sel_oi_one_hot_i[202] & i[175];
  assign _05075_ = sel_oi_one_hot_i[203] & i[191];
  assign _05076_ = _05075_ | _05074_;
  assign _05077_ = _05076_ | _05073_;
  assign _05078_ = sel_oi_one_hot_i[204] & i[207];
  assign _05079_ = sel_oi_one_hot_i[205] & i[223];
  assign _05080_ = _05079_ | _05078_;
  assign _05081_ = sel_oi_one_hot_i[206] & i[239];
  assign _05082_ = sel_oi_one_hot_i[207] & i[255];
  assign _05083_ = _05082_ | _05081_;
  assign _05084_ = _05083_ | _05080_;
  assign _05085_ = _05084_ | _05077_;
  assign o[207] = _05085_ | _05070_;
  assign _05086_ = sel_oi_one_hot_i[192] & i[14];
  assign _05087_ = sel_oi_one_hot_i[193] & i[30];
  assign _05088_ = _05087_ | _05086_;
  assign _05089_ = sel_oi_one_hot_i[194] & i[46];
  assign _05090_ = sel_oi_one_hot_i[195] & i[62];
  assign _05091_ = _05090_ | _05089_;
  assign _05092_ = _05091_ | _05088_;
  assign _05093_ = sel_oi_one_hot_i[196] & i[78];
  assign _05094_ = sel_oi_one_hot_i[197] & i[94];
  assign _05095_ = _05094_ | _05093_;
  assign _05096_ = sel_oi_one_hot_i[198] & i[110];
  assign _05097_ = sel_oi_one_hot_i[199] & i[126];
  assign _05098_ = _05097_ | _05096_;
  assign _05099_ = _05098_ | _05095_;
  assign _05100_ = _05099_ | _05092_;
  assign _05101_ = sel_oi_one_hot_i[200] & i[142];
  assign _05102_ = sel_oi_one_hot_i[201] & i[158];
  assign _05103_ = _05102_ | _05101_;
  assign _05104_ = sel_oi_one_hot_i[202] & i[174];
  assign _05105_ = sel_oi_one_hot_i[203] & i[190];
  assign _05106_ = _05105_ | _05104_;
  assign _05107_ = _05106_ | _05103_;
  assign _05108_ = sel_oi_one_hot_i[204] & i[206];
  assign _05109_ = sel_oi_one_hot_i[205] & i[222];
  assign _05110_ = _05109_ | _05108_;
  assign _05111_ = sel_oi_one_hot_i[206] & i[238];
  assign _05112_ = sel_oi_one_hot_i[207] & i[254];
  assign _05113_ = _05112_ | _05111_;
  assign _05114_ = _05113_ | _05110_;
  assign _05115_ = _05114_ | _05107_;
  assign o[206] = _05115_ | _05100_;
  assign _05116_ = i[15] & sel_oi_one_hot_i[16];
  assign _05117_ = i[31] & sel_oi_one_hot_i[17];
  assign _05118_ = _05117_ | _05116_;
  assign _05119_ = i[47] & sel_oi_one_hot_i[18];
  assign _05120_ = i[63] & sel_oi_one_hot_i[19];
  assign _05121_ = _05120_ | _05119_;
  assign _05122_ = _05121_ | _05118_;
  assign _05123_ = i[79] & sel_oi_one_hot_i[20];
  assign _05124_ = i[95] & sel_oi_one_hot_i[21];
  assign _05125_ = _05124_ | _05123_;
  assign _05126_ = i[111] & sel_oi_one_hot_i[22];
  assign _05127_ = i[127] & sel_oi_one_hot_i[23];
  assign _05128_ = _05127_ | _05126_;
  assign _05129_ = _05128_ | _05125_;
  assign _05130_ = _05129_ | _05122_;
  assign _05131_ = i[143] & sel_oi_one_hot_i[24];
  assign _05132_ = i[159] & sel_oi_one_hot_i[25];
  assign _05133_ = _05132_ | _05131_;
  assign _05134_ = i[175] & sel_oi_one_hot_i[26];
  assign _05135_ = i[191] & sel_oi_one_hot_i[27];
  assign _05136_ = _05135_ | _05134_;
  assign _05137_ = _05136_ | _05133_;
  assign _05138_ = i[207] & sel_oi_one_hot_i[28];
  assign _05139_ = i[223] & sel_oi_one_hot_i[29];
  assign _05140_ = _05139_ | _05138_;
  assign _05141_ = i[239] & sel_oi_one_hot_i[30];
  assign _05142_ = sel_oi_one_hot_i[31] & i[255];
  assign _05143_ = _05142_ | _05141_;
  assign _05144_ = _05143_ | _05140_;
  assign _05145_ = _05144_ | _05137_;
  assign o[31] = _05145_ | _05130_;
  assign _05146_ = sel_oi_one_hot_i[192] & i[13];
  assign _05147_ = sel_oi_one_hot_i[193] & i[29];
  assign _05148_ = _05147_ | _05146_;
  assign _05149_ = sel_oi_one_hot_i[194] & i[45];
  assign _05150_ = sel_oi_one_hot_i[195] & i[61];
  assign _05151_ = _05150_ | _05149_;
  assign _05152_ = _05151_ | _05148_;
  assign _05153_ = sel_oi_one_hot_i[196] & i[77];
  assign _05154_ = sel_oi_one_hot_i[197] & i[93];
  assign _05155_ = _05154_ | _05153_;
  assign _05156_ = sel_oi_one_hot_i[198] & i[109];
  assign _05157_ = sel_oi_one_hot_i[199] & i[125];
  assign _05158_ = _05157_ | _05156_;
  assign _05159_ = _05158_ | _05155_;
  assign _05160_ = _05159_ | _05152_;
  assign _05161_ = sel_oi_one_hot_i[200] & i[141];
  assign _05162_ = sel_oi_one_hot_i[201] & i[157];
  assign _05163_ = _05162_ | _05161_;
  assign _05164_ = sel_oi_one_hot_i[202] & i[173];
  assign _05165_ = sel_oi_one_hot_i[203] & i[189];
  assign _05166_ = _05165_ | _05164_;
  assign _05167_ = _05166_ | _05163_;
  assign _05168_ = sel_oi_one_hot_i[204] & i[205];
  assign _05169_ = sel_oi_one_hot_i[205] & i[221];
  assign _05170_ = _05169_ | _05168_;
  assign _05171_ = sel_oi_one_hot_i[206] & i[237];
  assign _05172_ = sel_oi_one_hot_i[207] & i[253];
  assign _05173_ = _05172_ | _05171_;
  assign _05174_ = _05173_ | _05170_;
  assign _05175_ = _05174_ | _05167_;
  assign o[205] = _05175_ | _05160_;
  assign _05176_ = sel_oi_one_hot_i[192] & i[12];
  assign _05177_ = sel_oi_one_hot_i[193] & i[28];
  assign _05178_ = _05177_ | _05176_;
  assign _05179_ = sel_oi_one_hot_i[194] & i[44];
  assign _05180_ = sel_oi_one_hot_i[195] & i[60];
  assign _05181_ = _05180_ | _05179_;
  assign _05182_ = _05181_ | _05178_;
  assign _05183_ = sel_oi_one_hot_i[196] & i[76];
  assign _05184_ = sel_oi_one_hot_i[197] & i[92];
  assign _05185_ = _05184_ | _05183_;
  assign _05186_ = sel_oi_one_hot_i[198] & i[108];
  assign _05187_ = sel_oi_one_hot_i[199] & i[124];
  assign _05188_ = _05187_ | _05186_;
  assign _05189_ = _05188_ | _05185_;
  assign _05190_ = _05189_ | _05182_;
  assign _05191_ = sel_oi_one_hot_i[200] & i[140];
  assign _05192_ = sel_oi_one_hot_i[201] & i[156];
  assign _05193_ = _05192_ | _05191_;
  assign _05194_ = sel_oi_one_hot_i[202] & i[172];
  assign _05195_ = sel_oi_one_hot_i[203] & i[188];
  assign _05196_ = _05195_ | _05194_;
  assign _05197_ = _05196_ | _05193_;
  assign _05198_ = sel_oi_one_hot_i[204] & i[204];
  assign _05199_ = sel_oi_one_hot_i[205] & i[220];
  assign _05200_ = _05199_ | _05198_;
  assign _05201_ = sel_oi_one_hot_i[206] & i[236];
  assign _05202_ = sel_oi_one_hot_i[207] & i[252];
  assign _05203_ = _05202_ | _05201_;
  assign _05204_ = _05203_ | _05200_;
  assign _05205_ = _05204_ | _05197_;
  assign o[204] = _05205_ | _05190_;
  assign _05206_ = sel_oi_one_hot_i[192] & i[11];
  assign _05207_ = sel_oi_one_hot_i[193] & i[27];
  assign _05208_ = _05207_ | _05206_;
  assign _05209_ = sel_oi_one_hot_i[194] & i[43];
  assign _05210_ = sel_oi_one_hot_i[195] & i[59];
  assign _05211_ = _05210_ | _05209_;
  assign _05212_ = _05211_ | _05208_;
  assign _05213_ = sel_oi_one_hot_i[196] & i[75];
  assign _05214_ = sel_oi_one_hot_i[197] & i[91];
  assign _05215_ = _05214_ | _05213_;
  assign _05216_ = sel_oi_one_hot_i[198] & i[107];
  assign _05217_ = sel_oi_one_hot_i[199] & i[123];
  assign _05218_ = _05217_ | _05216_;
  assign _05219_ = _05218_ | _05215_;
  assign _05220_ = _05219_ | _05212_;
  assign _05221_ = sel_oi_one_hot_i[200] & i[139];
  assign _05222_ = sel_oi_one_hot_i[201] & i[155];
  assign _05223_ = _05222_ | _05221_;
  assign _05224_ = sel_oi_one_hot_i[202] & i[171];
  assign _05225_ = sel_oi_one_hot_i[203] & i[187];
  assign _05226_ = _05225_ | _05224_;
  assign _05227_ = _05226_ | _05223_;
  assign _05228_ = sel_oi_one_hot_i[204] & i[203];
  assign _05229_ = sel_oi_one_hot_i[205] & i[219];
  assign _05230_ = _05229_ | _05228_;
  assign _05231_ = sel_oi_one_hot_i[206] & i[235];
  assign _05232_ = sel_oi_one_hot_i[207] & i[251];
  assign _05233_ = _05232_ | _05231_;
  assign _05234_ = _05233_ | _05230_;
  assign _05235_ = _05234_ | _05227_;
  assign o[203] = _05235_ | _05220_;
  assign _05236_ = sel_oi_one_hot_i[192] & i[10];
  assign _05237_ = sel_oi_one_hot_i[193] & i[26];
  assign _05238_ = _05237_ | _05236_;
  assign _05239_ = sel_oi_one_hot_i[194] & i[42];
  assign _05240_ = sel_oi_one_hot_i[195] & i[58];
  assign _05241_ = _05240_ | _05239_;
  assign _05242_ = _05241_ | _05238_;
  assign _05243_ = sel_oi_one_hot_i[196] & i[74];
  assign _05244_ = sel_oi_one_hot_i[197] & i[90];
  assign _05245_ = _05244_ | _05243_;
  assign _05246_ = sel_oi_one_hot_i[198] & i[106];
  assign _05247_ = sel_oi_one_hot_i[199] & i[122];
  assign _05248_ = _05247_ | _05246_;
  assign _05249_ = _05248_ | _05245_;
  assign _05250_ = _05249_ | _05242_;
  assign _05251_ = sel_oi_one_hot_i[200] & i[138];
  assign _05252_ = sel_oi_one_hot_i[201] & i[154];
  assign _05253_ = _05252_ | _05251_;
  assign _05254_ = sel_oi_one_hot_i[202] & i[170];
  assign _05255_ = sel_oi_one_hot_i[203] & i[186];
  assign _05256_ = _05255_ | _05254_;
  assign _05257_ = _05256_ | _05253_;
  assign _05258_ = sel_oi_one_hot_i[204] & i[202];
  assign _05259_ = sel_oi_one_hot_i[205] & i[218];
  assign _05260_ = _05259_ | _05258_;
  assign _05261_ = sel_oi_one_hot_i[206] & i[234];
  assign _05262_ = sel_oi_one_hot_i[207] & i[250];
  assign _05263_ = _05262_ | _05261_;
  assign _05264_ = _05263_ | _05260_;
  assign _05265_ = _05264_ | _05257_;
  assign o[202] = _05265_ | _05250_;
  assign _05266_ = sel_oi_one_hot_i[192] & i[9];
  assign _05267_ = sel_oi_one_hot_i[193] & i[25];
  assign _05268_ = _05267_ | _05266_;
  assign _05269_ = sel_oi_one_hot_i[194] & i[41];
  assign _05270_ = sel_oi_one_hot_i[195] & i[57];
  assign _05271_ = _05270_ | _05269_;
  assign _05272_ = _05271_ | _05268_;
  assign _05273_ = sel_oi_one_hot_i[196] & i[73];
  assign _05274_ = sel_oi_one_hot_i[197] & i[89];
  assign _05275_ = _05274_ | _05273_;
  assign _05276_ = sel_oi_one_hot_i[198] & i[105];
  assign _05277_ = sel_oi_one_hot_i[199] & i[121];
  assign _05278_ = _05277_ | _05276_;
  assign _05279_ = _05278_ | _05275_;
  assign _05280_ = _05279_ | _05272_;
  assign _05281_ = sel_oi_one_hot_i[200] & i[137];
  assign _05282_ = sel_oi_one_hot_i[201] & i[153];
  assign _05283_ = _05282_ | _05281_;
  assign _05284_ = sel_oi_one_hot_i[202] & i[169];
  assign _05285_ = sel_oi_one_hot_i[203] & i[185];
  assign _05286_ = _05285_ | _05284_;
  assign _05287_ = _05286_ | _05283_;
  assign _05288_ = sel_oi_one_hot_i[204] & i[201];
  assign _05289_ = sel_oi_one_hot_i[205] & i[217];
  assign _05290_ = _05289_ | _05288_;
  assign _05291_ = sel_oi_one_hot_i[206] & i[233];
  assign _05292_ = sel_oi_one_hot_i[207] & i[249];
  assign _05293_ = _05292_ | _05291_;
  assign _05294_ = _05293_ | _05290_;
  assign _05295_ = _05294_ | _05287_;
  assign o[201] = _05295_ | _05280_;
  assign _05296_ = sel_oi_one_hot_i[192] & i[8];
  assign _05297_ = sel_oi_one_hot_i[193] & i[24];
  assign _05298_ = _05297_ | _05296_;
  assign _05299_ = sel_oi_one_hot_i[194] & i[40];
  assign _05300_ = sel_oi_one_hot_i[195] & i[56];
  assign _05301_ = _05300_ | _05299_;
  assign _05302_ = _05301_ | _05298_;
  assign _05303_ = sel_oi_one_hot_i[196] & i[72];
  assign _05304_ = sel_oi_one_hot_i[197] & i[88];
  assign _05305_ = _05304_ | _05303_;
  assign _05306_ = sel_oi_one_hot_i[198] & i[104];
  assign _05307_ = sel_oi_one_hot_i[199] & i[120];
  assign _05308_ = _05307_ | _05306_;
  assign _05309_ = _05308_ | _05305_;
  assign _05310_ = _05309_ | _05302_;
  assign _05311_ = sel_oi_one_hot_i[200] & i[136];
  assign _05312_ = sel_oi_one_hot_i[201] & i[152];
  assign _05313_ = _05312_ | _05311_;
  assign _05314_ = sel_oi_one_hot_i[202] & i[168];
  assign _05315_ = sel_oi_one_hot_i[203] & i[184];
  assign _05316_ = _05315_ | _05314_;
  assign _05317_ = _05316_ | _05313_;
  assign _05318_ = sel_oi_one_hot_i[204] & i[200];
  assign _05319_ = sel_oi_one_hot_i[205] & i[216];
  assign _05320_ = _05319_ | _05318_;
  assign _05321_ = sel_oi_one_hot_i[206] & i[232];
  assign _05322_ = sel_oi_one_hot_i[207] & i[248];
  assign _05323_ = _05322_ | _05321_;
  assign _05324_ = _05323_ | _05320_;
  assign _05325_ = _05324_ | _05317_;
  assign o[200] = _05325_ | _05310_;
  assign _05326_ = sel_oi_one_hot_i[192] & i[7];
  assign _05327_ = sel_oi_one_hot_i[193] & i[23];
  assign _05328_ = _05327_ | _05326_;
  assign _05329_ = sel_oi_one_hot_i[194] & i[39];
  assign _05330_ = sel_oi_one_hot_i[195] & i[55];
  assign _05331_ = _05330_ | _05329_;
  assign _05332_ = _05331_ | _05328_;
  assign _05333_ = sel_oi_one_hot_i[196] & i[71];
  assign _05334_ = sel_oi_one_hot_i[197] & i[87];
  assign _05335_ = _05334_ | _05333_;
  assign _05336_ = sel_oi_one_hot_i[198] & i[103];
  assign _05337_ = sel_oi_one_hot_i[199] & i[119];
  assign _05338_ = _05337_ | _05336_;
  assign _05339_ = _05338_ | _05335_;
  assign _05340_ = _05339_ | _05332_;
  assign _05341_ = sel_oi_one_hot_i[200] & i[135];
  assign _05342_ = sel_oi_one_hot_i[201] & i[151];
  assign _05343_ = _05342_ | _05341_;
  assign _05344_ = sel_oi_one_hot_i[202] & i[167];
  assign _05345_ = sel_oi_one_hot_i[203] & i[183];
  assign _05346_ = _05345_ | _05344_;
  assign _05347_ = _05346_ | _05343_;
  assign _05348_ = sel_oi_one_hot_i[204] & i[199];
  assign _05349_ = sel_oi_one_hot_i[205] & i[215];
  assign _05350_ = _05349_ | _05348_;
  assign _05351_ = sel_oi_one_hot_i[206] & i[231];
  assign _05352_ = sel_oi_one_hot_i[207] & i[247];
  assign _05353_ = _05352_ | _05351_;
  assign _05354_ = _05353_ | _05350_;
  assign _05355_ = _05354_ | _05347_;
  assign o[199] = _05355_ | _05340_;
  assign _05356_ = sel_oi_one_hot_i[192] & i[6];
  assign _05357_ = sel_oi_one_hot_i[193] & i[22];
  assign _05358_ = _05357_ | _05356_;
  assign _05359_ = sel_oi_one_hot_i[194] & i[38];
  assign _05360_ = sel_oi_one_hot_i[195] & i[54];
  assign _05361_ = _05360_ | _05359_;
  assign _05362_ = _05361_ | _05358_;
  assign _05363_ = sel_oi_one_hot_i[196] & i[70];
  assign _05364_ = sel_oi_one_hot_i[197] & i[86];
  assign _05365_ = _05364_ | _05363_;
  assign _05366_ = sel_oi_one_hot_i[198] & i[102];
  assign _05367_ = sel_oi_one_hot_i[199] & i[118];
  assign _05368_ = _05367_ | _05366_;
  assign _05369_ = _05368_ | _05365_;
  assign _05370_ = _05369_ | _05362_;
  assign _05371_ = sel_oi_one_hot_i[200] & i[134];
  assign _05372_ = sel_oi_one_hot_i[201] & i[150];
  assign _05373_ = _05372_ | _05371_;
  assign _05374_ = sel_oi_one_hot_i[202] & i[166];
  assign _05375_ = sel_oi_one_hot_i[203] & i[182];
  assign _05376_ = _05375_ | _05374_;
  assign _05377_ = _05376_ | _05373_;
  assign _05378_ = sel_oi_one_hot_i[204] & i[198];
  assign _05379_ = sel_oi_one_hot_i[205] & i[214];
  assign _05380_ = _05379_ | _05378_;
  assign _05381_ = sel_oi_one_hot_i[206] & i[230];
  assign _05382_ = sel_oi_one_hot_i[207] & i[246];
  assign _05383_ = _05382_ | _05381_;
  assign _05384_ = _05383_ | _05380_;
  assign _05385_ = _05384_ | _05377_;
  assign o[198] = _05385_ | _05370_;
  assign _05386_ = sel_oi_one_hot_i[192] & i[5];
  assign _05387_ = sel_oi_one_hot_i[193] & i[21];
  assign _05388_ = _05387_ | _05386_;
  assign _05389_ = sel_oi_one_hot_i[194] & i[37];
  assign _05390_ = sel_oi_one_hot_i[195] & i[53];
  assign _05391_ = _05390_ | _05389_;
  assign _05392_ = _05391_ | _05388_;
  assign _05393_ = sel_oi_one_hot_i[196] & i[69];
  assign _05394_ = sel_oi_one_hot_i[197] & i[85];
  assign _05395_ = _05394_ | _05393_;
  assign _05396_ = sel_oi_one_hot_i[198] & i[101];
  assign _05397_ = sel_oi_one_hot_i[199] & i[117];
  assign _05398_ = _05397_ | _05396_;
  assign _05399_ = _05398_ | _05395_;
  assign _05400_ = _05399_ | _05392_;
  assign _05401_ = sel_oi_one_hot_i[200] & i[133];
  assign _05402_ = sel_oi_one_hot_i[201] & i[149];
  assign _05403_ = _05402_ | _05401_;
  assign _05404_ = sel_oi_one_hot_i[202] & i[165];
  assign _05405_ = sel_oi_one_hot_i[203] & i[181];
  assign _05406_ = _05405_ | _05404_;
  assign _05407_ = _05406_ | _05403_;
  assign _05408_ = sel_oi_one_hot_i[204] & i[197];
  assign _05409_ = sel_oi_one_hot_i[205] & i[213];
  assign _05410_ = _05409_ | _05408_;
  assign _05411_ = sel_oi_one_hot_i[206] & i[229];
  assign _05412_ = sel_oi_one_hot_i[207] & i[245];
  assign _05413_ = _05412_ | _05411_;
  assign _05414_ = _05413_ | _05410_;
  assign _05415_ = _05414_ | _05407_;
  assign o[197] = _05415_ | _05400_;
  assign _05416_ = sel_oi_one_hot_i[192] & i[4];
  assign _05417_ = sel_oi_one_hot_i[193] & i[20];
  assign _05418_ = _05417_ | _05416_;
  assign _05419_ = sel_oi_one_hot_i[194] & i[36];
  assign _05420_ = sel_oi_one_hot_i[195] & i[52];
  assign _05421_ = _05420_ | _05419_;
  assign _05422_ = _05421_ | _05418_;
  assign _05423_ = sel_oi_one_hot_i[196] & i[68];
  assign _05424_ = sel_oi_one_hot_i[197] & i[84];
  assign _05425_ = _05424_ | _05423_;
  assign _05426_ = sel_oi_one_hot_i[198] & i[100];
  assign _05427_ = sel_oi_one_hot_i[199] & i[116];
  assign _05428_ = _05427_ | _05426_;
  assign _05429_ = _05428_ | _05425_;
  assign _05430_ = _05429_ | _05422_;
  assign _05431_ = sel_oi_one_hot_i[200] & i[132];
  assign _05432_ = sel_oi_one_hot_i[201] & i[148];
  assign _05433_ = _05432_ | _05431_;
  assign _05434_ = sel_oi_one_hot_i[202] & i[164];
  assign _05435_ = sel_oi_one_hot_i[203] & i[180];
  assign _05436_ = _05435_ | _05434_;
  assign _05437_ = _05436_ | _05433_;
  assign _05438_ = sel_oi_one_hot_i[204] & i[196];
  assign _05439_ = sel_oi_one_hot_i[205] & i[212];
  assign _05440_ = _05439_ | _05438_;
  assign _05441_ = sel_oi_one_hot_i[206] & i[228];
  assign _05442_ = sel_oi_one_hot_i[207] & i[244];
  assign _05443_ = _05442_ | _05441_;
  assign _05444_ = _05443_ | _05440_;
  assign _05445_ = _05444_ | _05437_;
  assign o[196] = _05445_ | _05430_;
  assign _05446_ = i[14] & sel_oi_one_hot_i[16];
  assign _05447_ = i[30] & sel_oi_one_hot_i[17];
  assign _05448_ = _05447_ | _05446_;
  assign _05449_ = i[46] & sel_oi_one_hot_i[18];
  assign _05450_ = i[62] & sel_oi_one_hot_i[19];
  assign _05451_ = _05450_ | _05449_;
  assign _05452_ = _05451_ | _05448_;
  assign _05453_ = i[78] & sel_oi_one_hot_i[20];
  assign _05454_ = i[94] & sel_oi_one_hot_i[21];
  assign _05455_ = _05454_ | _05453_;
  assign _05456_ = i[110] & sel_oi_one_hot_i[22];
  assign _05457_ = i[126] & sel_oi_one_hot_i[23];
  assign _05458_ = _05457_ | _05456_;
  assign _05459_ = _05458_ | _05455_;
  assign _05460_ = _05459_ | _05452_;
  assign _05461_ = i[142] & sel_oi_one_hot_i[24];
  assign _05462_ = i[158] & sel_oi_one_hot_i[25];
  assign _05463_ = _05462_ | _05461_;
  assign _05464_ = i[174] & sel_oi_one_hot_i[26];
  assign _05465_ = i[190] & sel_oi_one_hot_i[27];
  assign _05466_ = _05465_ | _05464_;
  assign _05467_ = _05466_ | _05463_;
  assign _05468_ = i[206] & sel_oi_one_hot_i[28];
  assign _05469_ = i[222] & sel_oi_one_hot_i[29];
  assign _05470_ = _05469_ | _05468_;
  assign _05471_ = i[238] & sel_oi_one_hot_i[30];
  assign _05472_ = sel_oi_one_hot_i[31] & i[254];
  assign _05473_ = _05472_ | _05471_;
  assign _05474_ = _05473_ | _05470_;
  assign _05475_ = _05474_ | _05467_;
  assign o[30] = _05475_ | _05460_;
  assign _05476_ = sel_oi_one_hot_i[192] & i[3];
  assign _05477_ = sel_oi_one_hot_i[193] & i[19];
  assign _05478_ = _05477_ | _05476_;
  assign _05479_ = sel_oi_one_hot_i[194] & i[35];
  assign _05480_ = sel_oi_one_hot_i[195] & i[51];
  assign _05481_ = _05480_ | _05479_;
  assign _05482_ = _05481_ | _05478_;
  assign _05483_ = sel_oi_one_hot_i[196] & i[67];
  assign _05484_ = sel_oi_one_hot_i[197] & i[83];
  assign _05485_ = _05484_ | _05483_;
  assign _05486_ = sel_oi_one_hot_i[198] & i[99];
  assign _05487_ = sel_oi_one_hot_i[199] & i[115];
  assign _05488_ = _05487_ | _05486_;
  assign _05489_ = _05488_ | _05485_;
  assign _05490_ = _05489_ | _05482_;
  assign _05491_ = sel_oi_one_hot_i[200] & i[131];
  assign _05492_ = sel_oi_one_hot_i[201] & i[147];
  assign _05493_ = _05492_ | _05491_;
  assign _05494_ = sel_oi_one_hot_i[202] & i[163];
  assign _05495_ = sel_oi_one_hot_i[203] & i[179];
  assign _05496_ = _05495_ | _05494_;
  assign _05497_ = _05496_ | _05493_;
  assign _05498_ = sel_oi_one_hot_i[204] & i[195];
  assign _05499_ = sel_oi_one_hot_i[205] & i[211];
  assign _05500_ = _05499_ | _05498_;
  assign _05501_ = sel_oi_one_hot_i[206] & i[227];
  assign _05502_ = sel_oi_one_hot_i[207] & i[243];
  assign _05503_ = _05502_ | _05501_;
  assign _05504_ = _05503_ | _05500_;
  assign _05505_ = _05504_ | _05497_;
  assign o[195] = _05505_ | _05490_;
  assign _05506_ = sel_oi_one_hot_i[192] & i[2];
  assign _05507_ = sel_oi_one_hot_i[193] & i[18];
  assign _05508_ = _05507_ | _05506_;
  assign _05509_ = sel_oi_one_hot_i[194] & i[34];
  assign _05510_ = sel_oi_one_hot_i[195] & i[50];
  assign _05511_ = _05510_ | _05509_;
  assign _05512_ = _05511_ | _05508_;
  assign _05513_ = sel_oi_one_hot_i[196] & i[66];
  assign _05514_ = sel_oi_one_hot_i[197] & i[82];
  assign _05515_ = _05514_ | _05513_;
  assign _05516_ = sel_oi_one_hot_i[198] & i[98];
  assign _05517_ = sel_oi_one_hot_i[199] & i[114];
  assign _05518_ = _05517_ | _05516_;
  assign _05519_ = _05518_ | _05515_;
  assign _05520_ = _05519_ | _05512_;
  assign _05521_ = sel_oi_one_hot_i[200] & i[130];
  assign _05522_ = sel_oi_one_hot_i[201] & i[146];
  assign _05523_ = _05522_ | _05521_;
  assign _05524_ = sel_oi_one_hot_i[202] & i[162];
  assign _05525_ = sel_oi_one_hot_i[203] & i[178];
  assign _05526_ = _05525_ | _05524_;
  assign _05527_ = _05526_ | _05523_;
  assign _05528_ = sel_oi_one_hot_i[204] & i[194];
  assign _05529_ = sel_oi_one_hot_i[205] & i[210];
  assign _05530_ = _05529_ | _05528_;
  assign _05531_ = sel_oi_one_hot_i[206] & i[226];
  assign _05532_ = sel_oi_one_hot_i[207] & i[242];
  assign _05533_ = _05532_ | _05531_;
  assign _05534_ = _05533_ | _05530_;
  assign _05535_ = _05534_ | _05527_;
  assign o[194] = _05535_ | _05520_;
  assign _05536_ = sel_oi_one_hot_i[192] & i[1];
  assign _05537_ = sel_oi_one_hot_i[193] & i[17];
  assign _05538_ = _05537_ | _05536_;
  assign _05539_ = sel_oi_one_hot_i[194] & i[33];
  assign _05540_ = sel_oi_one_hot_i[195] & i[49];
  assign _05541_ = _05540_ | _05539_;
  assign _05542_ = _05541_ | _05538_;
  assign _05543_ = sel_oi_one_hot_i[196] & i[65];
  assign _05544_ = sel_oi_one_hot_i[197] & i[81];
  assign _05545_ = _05544_ | _05543_;
  assign _05546_ = sel_oi_one_hot_i[198] & i[97];
  assign _05547_ = sel_oi_one_hot_i[199] & i[113];
  assign _05548_ = _05547_ | _05546_;
  assign _05549_ = _05548_ | _05545_;
  assign _05550_ = _05549_ | _05542_;
  assign _05551_ = sel_oi_one_hot_i[200] & i[129];
  assign _05552_ = sel_oi_one_hot_i[201] & i[145];
  assign _05553_ = _05552_ | _05551_;
  assign _05554_ = sel_oi_one_hot_i[202] & i[161];
  assign _05555_ = sel_oi_one_hot_i[203] & i[177];
  assign _05556_ = _05555_ | _05554_;
  assign _05557_ = _05556_ | _05553_;
  assign _05558_ = sel_oi_one_hot_i[204] & i[193];
  assign _05559_ = sel_oi_one_hot_i[205] & i[209];
  assign _05560_ = _05559_ | _05558_;
  assign _05561_ = sel_oi_one_hot_i[206] & i[225];
  assign _05562_ = sel_oi_one_hot_i[207] & i[241];
  assign _05563_ = _05562_ | _05561_;
  assign _05564_ = _05563_ | _05560_;
  assign _05565_ = _05564_ | _05557_;
  assign o[193] = _05565_ | _05550_;
  assign _05566_ = sel_oi_one_hot_i[192] & i[0];
  assign _05567_ = sel_oi_one_hot_i[193] & i[16];
  assign _05568_ = _05567_ | _05566_;
  assign _05569_ = sel_oi_one_hot_i[194] & i[32];
  assign _05570_ = sel_oi_one_hot_i[195] & i[48];
  assign _05571_ = _05570_ | _05569_;
  assign _05572_ = _05571_ | _05568_;
  assign _05573_ = sel_oi_one_hot_i[196] & i[64];
  assign _05574_ = sel_oi_one_hot_i[197] & i[80];
  assign _05575_ = _05574_ | _05573_;
  assign _05576_ = sel_oi_one_hot_i[198] & i[96];
  assign _05577_ = sel_oi_one_hot_i[199] & i[112];
  assign _05578_ = _05577_ | _05576_;
  assign _05579_ = _05578_ | _05575_;
  assign _05580_ = _05579_ | _05572_;
  assign _05581_ = sel_oi_one_hot_i[200] & i[128];
  assign _05582_ = sel_oi_one_hot_i[201] & i[144];
  assign _05583_ = _05582_ | _05581_;
  assign _05584_ = sel_oi_one_hot_i[202] & i[160];
  assign _05585_ = sel_oi_one_hot_i[203] & i[176];
  assign _05586_ = _05585_ | _05584_;
  assign _05587_ = _05586_ | _05583_;
  assign _05588_ = sel_oi_one_hot_i[204] & i[192];
  assign _05589_ = sel_oi_one_hot_i[205] & i[208];
  assign _05590_ = _05589_ | _05588_;
  assign _05591_ = sel_oi_one_hot_i[206] & i[224];
  assign _05592_ = sel_oi_one_hot_i[207] & i[240];
  assign _05593_ = _05592_ | _05591_;
  assign _05594_ = _05593_ | _05590_;
  assign _05595_ = _05594_ | _05587_;
  assign o[192] = _05595_ | _05580_;
  assign _05596_ = i[13] & sel_oi_one_hot_i[16];
  assign _05597_ = i[29] & sel_oi_one_hot_i[17];
  assign _05598_ = _05597_ | _05596_;
  assign _05599_ = i[45] & sel_oi_one_hot_i[18];
  assign _05600_ = i[61] & sel_oi_one_hot_i[19];
  assign _05601_ = _05600_ | _05599_;
  assign _05602_ = _05601_ | _05598_;
  assign _05603_ = i[77] & sel_oi_one_hot_i[20];
  assign _05604_ = i[93] & sel_oi_one_hot_i[21];
  assign _05605_ = _05604_ | _05603_;
  assign _05606_ = i[109] & sel_oi_one_hot_i[22];
  assign _05607_ = i[125] & sel_oi_one_hot_i[23];
  assign _05608_ = _05607_ | _05606_;
  assign _05609_ = _05608_ | _05605_;
  assign _05610_ = _05609_ | _05602_;
  assign _05611_ = i[141] & sel_oi_one_hot_i[24];
  assign _05612_ = i[157] & sel_oi_one_hot_i[25];
  assign _05613_ = _05612_ | _05611_;
  assign _05614_ = i[173] & sel_oi_one_hot_i[26];
  assign _05615_ = i[189] & sel_oi_one_hot_i[27];
  assign _05616_ = _05615_ | _05614_;
  assign _05617_ = _05616_ | _05613_;
  assign _05618_ = i[205] & sel_oi_one_hot_i[28];
  assign _05619_ = i[221] & sel_oi_one_hot_i[29];
  assign _05620_ = _05619_ | _05618_;
  assign _05621_ = i[237] & sel_oi_one_hot_i[30];
  assign _05622_ = sel_oi_one_hot_i[31] & i[253];
  assign _05623_ = _05622_ | _05621_;
  assign _05624_ = _05623_ | _05620_;
  assign _05625_ = _05624_ | _05617_;
  assign o[29] = _05625_ | _05610_;
  assign _05626_ = sel_oi_one_hot_i[208] & i[15];
  assign _05627_ = sel_oi_one_hot_i[209] & i[31];
  assign _05628_ = _05627_ | _05626_;
  assign _05629_ = sel_oi_one_hot_i[210] & i[47];
  assign _05630_ = sel_oi_one_hot_i[211] & i[63];
  assign _05631_ = _05630_ | _05629_;
  assign _05632_ = _05631_ | _05628_;
  assign _05633_ = sel_oi_one_hot_i[212] & i[79];
  assign _05634_ = sel_oi_one_hot_i[213] & i[95];
  assign _05635_ = _05634_ | _05633_;
  assign _05636_ = sel_oi_one_hot_i[214] & i[111];
  assign _05637_ = sel_oi_one_hot_i[215] & i[127];
  assign _05638_ = _05637_ | _05636_;
  assign _05639_ = _05638_ | _05635_;
  assign _05640_ = _05639_ | _05632_;
  assign _05641_ = sel_oi_one_hot_i[216] & i[143];
  assign _05642_ = sel_oi_one_hot_i[217] & i[159];
  assign _05643_ = _05642_ | _05641_;
  assign _05644_ = sel_oi_one_hot_i[218] & i[175];
  assign _05645_ = sel_oi_one_hot_i[219] & i[191];
  assign _05646_ = _05645_ | _05644_;
  assign _05647_ = _05646_ | _05643_;
  assign _05648_ = sel_oi_one_hot_i[220] & i[207];
  assign _05649_ = sel_oi_one_hot_i[221] & i[223];
  assign _05650_ = _05649_ | _05648_;
  assign _05651_ = sel_oi_one_hot_i[222] & i[239];
  assign _05652_ = sel_oi_one_hot_i[223] & i[255];
  assign _05653_ = _05652_ | _05651_;
  assign _05654_ = _05653_ | _05650_;
  assign _05655_ = _05654_ | _05647_;
  assign o[223] = _05655_ | _05640_;
  assign _05656_ = sel_oi_one_hot_i[208] & i[14];
  assign _05657_ = sel_oi_one_hot_i[209] & i[30];
  assign _05658_ = _05657_ | _05656_;
  assign _05659_ = sel_oi_one_hot_i[210] & i[46];
  assign _05660_ = sel_oi_one_hot_i[211] & i[62];
  assign _05661_ = _05660_ | _05659_;
  assign _05662_ = _05661_ | _05658_;
  assign _05663_ = sel_oi_one_hot_i[212] & i[78];
  assign _05664_ = sel_oi_one_hot_i[213] & i[94];
  assign _05665_ = _05664_ | _05663_;
  assign _05666_ = sel_oi_one_hot_i[214] & i[110];
  assign _05667_ = sel_oi_one_hot_i[215] & i[126];
  assign _05668_ = _05667_ | _05666_;
  assign _05669_ = _05668_ | _05665_;
  assign _05670_ = _05669_ | _05662_;
  assign _05671_ = sel_oi_one_hot_i[216] & i[142];
  assign _05672_ = sel_oi_one_hot_i[217] & i[158];
  assign _05673_ = _05672_ | _05671_;
  assign _05674_ = sel_oi_one_hot_i[218] & i[174];
  assign _05675_ = sel_oi_one_hot_i[219] & i[190];
  assign _05676_ = _05675_ | _05674_;
  assign _05677_ = _05676_ | _05673_;
  assign _05678_ = sel_oi_one_hot_i[220] & i[206];
  assign _05679_ = sel_oi_one_hot_i[221] & i[222];
  assign _05680_ = _05679_ | _05678_;
  assign _05681_ = sel_oi_one_hot_i[222] & i[238];
  assign _05682_ = sel_oi_one_hot_i[223] & i[254];
  assign _05683_ = _05682_ | _05681_;
  assign _05684_ = _05683_ | _05680_;
  assign _05685_ = _05684_ | _05677_;
  assign o[222] = _05685_ | _05670_;
  assign _05686_ = sel_oi_one_hot_i[208] & i[13];
  assign _05687_ = sel_oi_one_hot_i[209] & i[29];
  assign _05688_ = _05687_ | _05686_;
  assign _05689_ = sel_oi_one_hot_i[210] & i[45];
  assign _05690_ = sel_oi_one_hot_i[211] & i[61];
  assign _05691_ = _05690_ | _05689_;
  assign _05692_ = _05691_ | _05688_;
  assign _05693_ = sel_oi_one_hot_i[212] & i[77];
  assign _05694_ = sel_oi_one_hot_i[213] & i[93];
  assign _05695_ = _05694_ | _05693_;
  assign _05696_ = sel_oi_one_hot_i[214] & i[109];
  assign _05697_ = sel_oi_one_hot_i[215] & i[125];
  assign _05698_ = _05697_ | _05696_;
  assign _05699_ = _05698_ | _05695_;
  assign _05700_ = _05699_ | _05692_;
  assign _05701_ = sel_oi_one_hot_i[216] & i[141];
  assign _05702_ = sel_oi_one_hot_i[217] & i[157];
  assign _05703_ = _05702_ | _05701_;
  assign _05704_ = sel_oi_one_hot_i[218] & i[173];
  assign _05705_ = sel_oi_one_hot_i[219] & i[189];
  assign _05706_ = _05705_ | _05704_;
  assign _05707_ = _05706_ | _05703_;
  assign _05708_ = sel_oi_one_hot_i[220] & i[205];
  assign _05709_ = sel_oi_one_hot_i[221] & i[221];
  assign _05710_ = _05709_ | _05708_;
  assign _05711_ = sel_oi_one_hot_i[222] & i[237];
  assign _05712_ = sel_oi_one_hot_i[223] & i[253];
  assign _05713_ = _05712_ | _05711_;
  assign _05714_ = _05713_ | _05710_;
  assign _05715_ = _05714_ | _05707_;
  assign o[221] = _05715_ | _05700_;
  assign _05716_ = i[12] & sel_oi_one_hot_i[16];
  assign _05717_ = i[28] & sel_oi_one_hot_i[17];
  assign _05718_ = _05717_ | _05716_;
  assign _05719_ = i[44] & sel_oi_one_hot_i[18];
  assign _05720_ = i[60] & sel_oi_one_hot_i[19];
  assign _05721_ = _05720_ | _05719_;
  assign _05722_ = _05721_ | _05718_;
  assign _05723_ = i[76] & sel_oi_one_hot_i[20];
  assign _05724_ = i[92] & sel_oi_one_hot_i[21];
  assign _05725_ = _05724_ | _05723_;
  assign _05726_ = i[108] & sel_oi_one_hot_i[22];
  assign _05727_ = i[124] & sel_oi_one_hot_i[23];
  assign _05728_ = _05727_ | _05726_;
  assign _05729_ = _05728_ | _05725_;
  assign _05730_ = _05729_ | _05722_;
  assign _05731_ = i[140] & sel_oi_one_hot_i[24];
  assign _05732_ = i[156] & sel_oi_one_hot_i[25];
  assign _05733_ = _05732_ | _05731_;
  assign _05734_ = i[172] & sel_oi_one_hot_i[26];
  assign _05735_ = i[188] & sel_oi_one_hot_i[27];
  assign _05736_ = _05735_ | _05734_;
  assign _05737_ = _05736_ | _05733_;
  assign _05738_ = i[204] & sel_oi_one_hot_i[28];
  assign _05739_ = i[220] & sel_oi_one_hot_i[29];
  assign _05740_ = _05739_ | _05738_;
  assign _05741_ = i[236] & sel_oi_one_hot_i[30];
  assign _05742_ = sel_oi_one_hot_i[31] & i[252];
  assign _05743_ = _05742_ | _05741_;
  assign _05744_ = _05743_ | _05740_;
  assign _05745_ = _05744_ | _05737_;
  assign o[28] = _05745_ | _05730_;
  assign _05746_ = sel_oi_one_hot_i[208] & i[12];
  assign _05747_ = sel_oi_one_hot_i[209] & i[28];
  assign _05748_ = _05747_ | _05746_;
  assign _05749_ = sel_oi_one_hot_i[210] & i[44];
  assign _05750_ = sel_oi_one_hot_i[211] & i[60];
  assign _05751_ = _05750_ | _05749_;
  assign _05752_ = _05751_ | _05748_;
  assign _05753_ = sel_oi_one_hot_i[212] & i[76];
  assign _05754_ = sel_oi_one_hot_i[213] & i[92];
  assign _05755_ = _05754_ | _05753_;
  assign _05756_ = sel_oi_one_hot_i[214] & i[108];
  assign _05757_ = sel_oi_one_hot_i[215] & i[124];
  assign _05758_ = _05757_ | _05756_;
  assign _05759_ = _05758_ | _05755_;
  assign _05760_ = _05759_ | _05752_;
  assign _05761_ = sel_oi_one_hot_i[216] & i[140];
  assign _05762_ = sel_oi_one_hot_i[217] & i[156];
  assign _05763_ = _05762_ | _05761_;
  assign _05764_ = sel_oi_one_hot_i[218] & i[172];
  assign _05765_ = sel_oi_one_hot_i[219] & i[188];
  assign _05766_ = _05765_ | _05764_;
  assign _05767_ = _05766_ | _05763_;
  assign _05768_ = sel_oi_one_hot_i[220] & i[204];
  assign _05769_ = sel_oi_one_hot_i[221] & i[220];
  assign _05770_ = _05769_ | _05768_;
  assign _05771_ = sel_oi_one_hot_i[222] & i[236];
  assign _05772_ = sel_oi_one_hot_i[223] & i[252];
  assign _05773_ = _05772_ | _05771_;
  assign _05774_ = _05773_ | _05770_;
  assign _05775_ = _05774_ | _05767_;
  assign o[220] = _05775_ | _05760_;
  assign _05776_ = sel_oi_one_hot_i[208] & i[11];
  assign _05777_ = sel_oi_one_hot_i[209] & i[27];
  assign _05778_ = _05777_ | _05776_;
  assign _05779_ = sel_oi_one_hot_i[210] & i[43];
  assign _05780_ = sel_oi_one_hot_i[211] & i[59];
  assign _05781_ = _05780_ | _05779_;
  assign _05782_ = _05781_ | _05778_;
  assign _05783_ = sel_oi_one_hot_i[212] & i[75];
  assign _05784_ = sel_oi_one_hot_i[213] & i[91];
  assign _05785_ = _05784_ | _05783_;
  assign _05786_ = sel_oi_one_hot_i[214] & i[107];
  assign _05787_ = sel_oi_one_hot_i[215] & i[123];
  assign _05788_ = _05787_ | _05786_;
  assign _05789_ = _05788_ | _05785_;
  assign _05790_ = _05789_ | _05782_;
  assign _05791_ = sel_oi_one_hot_i[216] & i[139];
  assign _05792_ = sel_oi_one_hot_i[217] & i[155];
  assign _05793_ = _05792_ | _05791_;
  assign _05794_ = sel_oi_one_hot_i[218] & i[171];
  assign _05795_ = sel_oi_one_hot_i[219] & i[187];
  assign _05796_ = _05795_ | _05794_;
  assign _05797_ = _05796_ | _05793_;
  assign _05798_ = sel_oi_one_hot_i[220] & i[203];
  assign _05799_ = sel_oi_one_hot_i[221] & i[219];
  assign _05800_ = _05799_ | _05798_;
  assign _05801_ = sel_oi_one_hot_i[222] & i[235];
  assign _05802_ = sel_oi_one_hot_i[223] & i[251];
  assign _05803_ = _05802_ | _05801_;
  assign _05804_ = _05803_ | _05800_;
  assign _05805_ = _05804_ | _05797_;
  assign o[219] = _05805_ | _05790_;
  assign _05806_ = sel_oi_one_hot_i[208] & i[10];
  assign _05807_ = sel_oi_one_hot_i[209] & i[26];
  assign _05808_ = _05807_ | _05806_;
  assign _05809_ = sel_oi_one_hot_i[210] & i[42];
  assign _05810_ = sel_oi_one_hot_i[211] & i[58];
  assign _05811_ = _05810_ | _05809_;
  assign _05812_ = _05811_ | _05808_;
  assign _05813_ = sel_oi_one_hot_i[212] & i[74];
  assign _05814_ = sel_oi_one_hot_i[213] & i[90];
  assign _05815_ = _05814_ | _05813_;
  assign _05816_ = sel_oi_one_hot_i[214] & i[106];
  assign _05817_ = sel_oi_one_hot_i[215] & i[122];
  assign _05818_ = _05817_ | _05816_;
  assign _05819_ = _05818_ | _05815_;
  assign _05820_ = _05819_ | _05812_;
  assign _05821_ = sel_oi_one_hot_i[216] & i[138];
  assign _05822_ = sel_oi_one_hot_i[217] & i[154];
  assign _05823_ = _05822_ | _05821_;
  assign _05824_ = sel_oi_one_hot_i[218] & i[170];
  assign _05825_ = sel_oi_one_hot_i[219] & i[186];
  assign _05826_ = _05825_ | _05824_;
  assign _05827_ = _05826_ | _05823_;
  assign _05828_ = sel_oi_one_hot_i[220] & i[202];
  assign _05829_ = sel_oi_one_hot_i[221] & i[218];
  assign _05830_ = _05829_ | _05828_;
  assign _05831_ = sel_oi_one_hot_i[222] & i[234];
  assign _05832_ = sel_oi_one_hot_i[223] & i[250];
  assign _05833_ = _05832_ | _05831_;
  assign _05834_ = _05833_ | _05830_;
  assign _05835_ = _05834_ | _05827_;
  assign o[218] = _05835_ | _05820_;
  assign _05836_ = sel_oi_one_hot_i[208] & i[9];
  assign _05837_ = sel_oi_one_hot_i[209] & i[25];
  assign _05838_ = _05837_ | _05836_;
  assign _05839_ = sel_oi_one_hot_i[210] & i[41];
  assign _05840_ = sel_oi_one_hot_i[211] & i[57];
  assign _05841_ = _05840_ | _05839_;
  assign _05842_ = _05841_ | _05838_;
  assign _05843_ = sel_oi_one_hot_i[212] & i[73];
  assign _05844_ = sel_oi_one_hot_i[213] & i[89];
  assign _05845_ = _05844_ | _05843_;
  assign _05846_ = sel_oi_one_hot_i[214] & i[105];
  assign _05847_ = sel_oi_one_hot_i[215] & i[121];
  assign _05848_ = _05847_ | _05846_;
  assign _05849_ = _05848_ | _05845_;
  assign _05850_ = _05849_ | _05842_;
  assign _05851_ = sel_oi_one_hot_i[216] & i[137];
  assign _05852_ = sel_oi_one_hot_i[217] & i[153];
  assign _05853_ = _05852_ | _05851_;
  assign _05854_ = sel_oi_one_hot_i[218] & i[169];
  assign _05855_ = sel_oi_one_hot_i[219] & i[185];
  assign _05856_ = _05855_ | _05854_;
  assign _05857_ = _05856_ | _05853_;
  assign _05858_ = sel_oi_one_hot_i[220] & i[201];
  assign _05859_ = sel_oi_one_hot_i[221] & i[217];
  assign _05860_ = _05859_ | _05858_;
  assign _05861_ = sel_oi_one_hot_i[222] & i[233];
  assign _05862_ = sel_oi_one_hot_i[223] & i[249];
  assign _05863_ = _05862_ | _05861_;
  assign _05864_ = _05863_ | _05860_;
  assign _05865_ = _05864_ | _05857_;
  assign o[217] = _05865_ | _05850_;
  assign _05866_ = sel_oi_one_hot_i[208] & i[8];
  assign _05867_ = sel_oi_one_hot_i[209] & i[24];
  assign _05868_ = _05867_ | _05866_;
  assign _05869_ = sel_oi_one_hot_i[210] & i[40];
  assign _05870_ = sel_oi_one_hot_i[211] & i[56];
  assign _05871_ = _05870_ | _05869_;
  assign _05872_ = _05871_ | _05868_;
  assign _05873_ = sel_oi_one_hot_i[212] & i[72];
  assign _05874_ = sel_oi_one_hot_i[213] & i[88];
  assign _05875_ = _05874_ | _05873_;
  assign _05876_ = sel_oi_one_hot_i[214] & i[104];
  assign _05877_ = sel_oi_one_hot_i[215] & i[120];
  assign _05878_ = _05877_ | _05876_;
  assign _05879_ = _05878_ | _05875_;
  assign _05880_ = _05879_ | _05872_;
  assign _05881_ = sel_oi_one_hot_i[216] & i[136];
  assign _05882_ = sel_oi_one_hot_i[217] & i[152];
  assign _05883_ = _05882_ | _05881_;
  assign _05884_ = sel_oi_one_hot_i[218] & i[168];
  assign _05885_ = sel_oi_one_hot_i[219] & i[184];
  assign _05886_ = _05885_ | _05884_;
  assign _05887_ = _05886_ | _05883_;
  assign _05888_ = sel_oi_one_hot_i[220] & i[200];
  assign _05889_ = sel_oi_one_hot_i[221] & i[216];
  assign _05890_ = _05889_ | _05888_;
  assign _05891_ = sel_oi_one_hot_i[222] & i[232];
  assign _05892_ = sel_oi_one_hot_i[223] & i[248];
  assign _05893_ = _05892_ | _05891_;
  assign _05894_ = _05893_ | _05890_;
  assign _05895_ = _05894_ | _05887_;
  assign o[216] = _05895_ | _05880_;
  assign _05896_ = sel_oi_one_hot_i[208] & i[7];
  assign _05897_ = sel_oi_one_hot_i[209] & i[23];
  assign _05898_ = _05897_ | _05896_;
  assign _05899_ = sel_oi_one_hot_i[210] & i[39];
  assign _05900_ = sel_oi_one_hot_i[211] & i[55];
  assign _05901_ = _05900_ | _05899_;
  assign _05902_ = _05901_ | _05898_;
  assign _05903_ = sel_oi_one_hot_i[212] & i[71];
  assign _05904_ = sel_oi_one_hot_i[213] & i[87];
  assign _05905_ = _05904_ | _05903_;
  assign _05906_ = sel_oi_one_hot_i[214] & i[103];
  assign _05907_ = sel_oi_one_hot_i[215] & i[119];
  assign _05908_ = _05907_ | _05906_;
  assign _05909_ = _05908_ | _05905_;
  assign _05910_ = _05909_ | _05902_;
  assign _05911_ = sel_oi_one_hot_i[216] & i[135];
  assign _05912_ = sel_oi_one_hot_i[217] & i[151];
  assign _05913_ = _05912_ | _05911_;
  assign _05914_ = sel_oi_one_hot_i[218] & i[167];
  assign _05915_ = sel_oi_one_hot_i[219] & i[183];
  assign _05916_ = _05915_ | _05914_;
  assign _05917_ = _05916_ | _05913_;
  assign _05918_ = sel_oi_one_hot_i[220] & i[199];
  assign _05919_ = sel_oi_one_hot_i[221] & i[215];
  assign _05920_ = _05919_ | _05918_;
  assign _05921_ = sel_oi_one_hot_i[222] & i[231];
  assign _05922_ = sel_oi_one_hot_i[223] & i[247];
  assign _05923_ = _05922_ | _05921_;
  assign _05924_ = _05923_ | _05920_;
  assign _05925_ = _05924_ | _05917_;
  assign o[215] = _05925_ | _05910_;
  assign _05926_ = sel_oi_one_hot_i[208] & i[6];
  assign _05927_ = sel_oi_one_hot_i[209] & i[22];
  assign _05928_ = _05927_ | _05926_;
  assign _05929_ = sel_oi_one_hot_i[210] & i[38];
  assign _05930_ = sel_oi_one_hot_i[211] & i[54];
  assign _05931_ = _05930_ | _05929_;
  assign _05932_ = _05931_ | _05928_;
  assign _05933_ = sel_oi_one_hot_i[212] & i[70];
  assign _05934_ = sel_oi_one_hot_i[213] & i[86];
  assign _05935_ = _05934_ | _05933_;
  assign _05936_ = sel_oi_one_hot_i[214] & i[102];
  assign _05937_ = sel_oi_one_hot_i[215] & i[118];
  assign _05938_ = _05937_ | _05936_;
  assign _05939_ = _05938_ | _05935_;
  assign _05940_ = _05939_ | _05932_;
  assign _05941_ = sel_oi_one_hot_i[216] & i[134];
  assign _05942_ = sel_oi_one_hot_i[217] & i[150];
  assign _05943_ = _05942_ | _05941_;
  assign _05944_ = sel_oi_one_hot_i[218] & i[166];
  assign _05945_ = sel_oi_one_hot_i[219] & i[182];
  assign _05946_ = _05945_ | _05944_;
  assign _05947_ = _05946_ | _05943_;
  assign _05948_ = sel_oi_one_hot_i[220] & i[198];
  assign _05949_ = sel_oi_one_hot_i[221] & i[214];
  assign _05950_ = _05949_ | _05948_;
  assign _05951_ = sel_oi_one_hot_i[222] & i[230];
  assign _05952_ = sel_oi_one_hot_i[223] & i[246];
  assign _05953_ = _05952_ | _05951_;
  assign _05954_ = _05953_ | _05950_;
  assign _05955_ = _05954_ | _05947_;
  assign o[214] = _05955_ | _05940_;
  assign _05956_ = sel_oi_one_hot_i[208] & i[5];
  assign _05957_ = sel_oi_one_hot_i[209] & i[21];
  assign _05958_ = _05957_ | _05956_;
  assign _05959_ = sel_oi_one_hot_i[210] & i[37];
  assign _05960_ = sel_oi_one_hot_i[211] & i[53];
  assign _05961_ = _05960_ | _05959_;
  assign _05962_ = _05961_ | _05958_;
  assign _05963_ = sel_oi_one_hot_i[212] & i[69];
  assign _05964_ = sel_oi_one_hot_i[213] & i[85];
  assign _05965_ = _05964_ | _05963_;
  assign _05966_ = sel_oi_one_hot_i[214] & i[101];
  assign _05967_ = sel_oi_one_hot_i[215] & i[117];
  assign _05968_ = _05967_ | _05966_;
  assign _05969_ = _05968_ | _05965_;
  assign _05970_ = _05969_ | _05962_;
  assign _05971_ = sel_oi_one_hot_i[216] & i[133];
  assign _05972_ = sel_oi_one_hot_i[217] & i[149];
  assign _05973_ = _05972_ | _05971_;
  assign _05974_ = sel_oi_one_hot_i[218] & i[165];
  assign _05975_ = sel_oi_one_hot_i[219] & i[181];
  assign _05976_ = _05975_ | _05974_;
  assign _05977_ = _05976_ | _05973_;
  assign _05978_ = sel_oi_one_hot_i[220] & i[197];
  assign _05979_ = sel_oi_one_hot_i[221] & i[213];
  assign _05980_ = _05979_ | _05978_;
  assign _05981_ = sel_oi_one_hot_i[222] & i[229];
  assign _05982_ = sel_oi_one_hot_i[223] & i[245];
  assign _05983_ = _05982_ | _05981_;
  assign _05984_ = _05983_ | _05980_;
  assign _05985_ = _05984_ | _05977_;
  assign o[213] = _05985_ | _05970_;
  assign _05986_ = sel_oi_one_hot_i[208] & i[4];
  assign _05987_ = sel_oi_one_hot_i[209] & i[20];
  assign _05988_ = _05987_ | _05986_;
  assign _05989_ = sel_oi_one_hot_i[210] & i[36];
  assign _05990_ = sel_oi_one_hot_i[211] & i[52];
  assign _05991_ = _05990_ | _05989_;
  assign _05992_ = _05991_ | _05988_;
  assign _05993_ = sel_oi_one_hot_i[212] & i[68];
  assign _05994_ = sel_oi_one_hot_i[213] & i[84];
  assign _05995_ = _05994_ | _05993_;
  assign _05996_ = sel_oi_one_hot_i[214] & i[100];
  assign _05997_ = sel_oi_one_hot_i[215] & i[116];
  assign _05998_ = _05997_ | _05996_;
  assign _05999_ = _05998_ | _05995_;
  assign _06000_ = _05999_ | _05992_;
  assign _06001_ = sel_oi_one_hot_i[216] & i[132];
  assign _06002_ = sel_oi_one_hot_i[217] & i[148];
  assign _06003_ = _06002_ | _06001_;
  assign _06004_ = sel_oi_one_hot_i[218] & i[164];
  assign _06005_ = sel_oi_one_hot_i[219] & i[180];
  assign _06006_ = _06005_ | _06004_;
  assign _06007_ = _06006_ | _06003_;
  assign _06008_ = sel_oi_one_hot_i[220] & i[196];
  assign _06009_ = sel_oi_one_hot_i[221] & i[212];
  assign _06010_ = _06009_ | _06008_;
  assign _06011_ = sel_oi_one_hot_i[222] & i[228];
  assign _06012_ = sel_oi_one_hot_i[223] & i[244];
  assign _06013_ = _06012_ | _06011_;
  assign _06014_ = _06013_ | _06010_;
  assign _06015_ = _06014_ | _06007_;
  assign o[212] = _06015_ | _06000_;
  assign _06016_ = sel_oi_one_hot_i[208] & i[3];
  assign _06017_ = sel_oi_one_hot_i[209] & i[19];
  assign _06018_ = _06017_ | _06016_;
  assign _06019_ = sel_oi_one_hot_i[210] & i[35];
  assign _06020_ = sel_oi_one_hot_i[211] & i[51];
  assign _06021_ = _06020_ | _06019_;
  assign _06022_ = _06021_ | _06018_;
  assign _06023_ = sel_oi_one_hot_i[212] & i[67];
  assign _06024_ = sel_oi_one_hot_i[213] & i[83];
  assign _06025_ = _06024_ | _06023_;
  assign _06026_ = sel_oi_one_hot_i[214] & i[99];
  assign _06027_ = sel_oi_one_hot_i[215] & i[115];
  assign _06028_ = _06027_ | _06026_;
  assign _06029_ = _06028_ | _06025_;
  assign _06030_ = _06029_ | _06022_;
  assign _06031_ = sel_oi_one_hot_i[216] & i[131];
  assign _06032_ = sel_oi_one_hot_i[217] & i[147];
  assign _06033_ = _06032_ | _06031_;
  assign _06034_ = sel_oi_one_hot_i[218] & i[163];
  assign _06035_ = sel_oi_one_hot_i[219] & i[179];
  assign _06036_ = _06035_ | _06034_;
  assign _06037_ = _06036_ | _06033_;
  assign _06038_ = sel_oi_one_hot_i[220] & i[195];
  assign _06039_ = sel_oi_one_hot_i[221] & i[211];
  assign _06040_ = _06039_ | _06038_;
  assign _06041_ = sel_oi_one_hot_i[222] & i[227];
  assign _06042_ = sel_oi_one_hot_i[223] & i[243];
  assign _06043_ = _06042_ | _06041_;
  assign _06044_ = _06043_ | _06040_;
  assign _06045_ = _06044_ | _06037_;
  assign o[211] = _06045_ | _06030_;
  assign _06046_ = i[11] & sel_oi_one_hot_i[16];
  assign _06047_ = i[27] & sel_oi_one_hot_i[17];
  assign _06048_ = _06047_ | _06046_;
  assign _06049_ = i[43] & sel_oi_one_hot_i[18];
  assign _06050_ = i[59] & sel_oi_one_hot_i[19];
  assign _06051_ = _06050_ | _06049_;
  assign _06052_ = _06051_ | _06048_;
  assign _06053_ = i[75] & sel_oi_one_hot_i[20];
  assign _06054_ = i[91] & sel_oi_one_hot_i[21];
  assign _06055_ = _06054_ | _06053_;
  assign _06056_ = i[107] & sel_oi_one_hot_i[22];
  assign _06057_ = i[123] & sel_oi_one_hot_i[23];
  assign _06058_ = _06057_ | _06056_;
  assign _06059_ = _06058_ | _06055_;
  assign _06060_ = _06059_ | _06052_;
  assign _06061_ = i[139] & sel_oi_one_hot_i[24];
  assign _06062_ = i[155] & sel_oi_one_hot_i[25];
  assign _06063_ = _06062_ | _06061_;
  assign _06064_ = i[171] & sel_oi_one_hot_i[26];
  assign _06065_ = i[187] & sel_oi_one_hot_i[27];
  assign _06066_ = _06065_ | _06064_;
  assign _06067_ = _06066_ | _06063_;
  assign _06068_ = i[203] & sel_oi_one_hot_i[28];
  assign _06069_ = i[219] & sel_oi_one_hot_i[29];
  assign _06070_ = _06069_ | _06068_;
  assign _06071_ = i[235] & sel_oi_one_hot_i[30];
  assign _06072_ = sel_oi_one_hot_i[31] & i[251];
  assign _06073_ = _06072_ | _06071_;
  assign _06074_ = _06073_ | _06070_;
  assign _06075_ = _06074_ | _06067_;
  assign o[27] = _06075_ | _06060_;
  assign _06076_ = sel_oi_one_hot_i[208] & i[2];
  assign _06077_ = sel_oi_one_hot_i[209] & i[18];
  assign _06078_ = _06077_ | _06076_;
  assign _06079_ = sel_oi_one_hot_i[210] & i[34];
  assign _06080_ = sel_oi_one_hot_i[211] & i[50];
  assign _06081_ = _06080_ | _06079_;
  assign _06082_ = _06081_ | _06078_;
  assign _06083_ = sel_oi_one_hot_i[212] & i[66];
  assign _06084_ = sel_oi_one_hot_i[213] & i[82];
  assign _06085_ = _06084_ | _06083_;
  assign _06086_ = sel_oi_one_hot_i[214] & i[98];
  assign _06087_ = sel_oi_one_hot_i[215] & i[114];
  assign _06088_ = _06087_ | _06086_;
  assign _06089_ = _06088_ | _06085_;
  assign _06090_ = _06089_ | _06082_;
  assign _06091_ = sel_oi_one_hot_i[216] & i[130];
  assign _06092_ = sel_oi_one_hot_i[217] & i[146];
  assign _06093_ = _06092_ | _06091_;
  assign _06094_ = sel_oi_one_hot_i[218] & i[162];
  assign _06095_ = sel_oi_one_hot_i[219] & i[178];
  assign _06096_ = _06095_ | _06094_;
  assign _06097_ = _06096_ | _06093_;
  assign _06098_ = sel_oi_one_hot_i[220] & i[194];
  assign _06099_ = sel_oi_one_hot_i[221] & i[210];
  assign _06100_ = _06099_ | _06098_;
  assign _06101_ = sel_oi_one_hot_i[222] & i[226];
  assign _06102_ = sel_oi_one_hot_i[223] & i[242];
  assign _06103_ = _06102_ | _06101_;
  assign _06104_ = _06103_ | _06100_;
  assign _06105_ = _06104_ | _06097_;
  assign o[210] = _06105_ | _06090_;
  assign _06106_ = sel_oi_one_hot_i[208] & i[1];
  assign _06107_ = sel_oi_one_hot_i[209] & i[17];
  assign _06108_ = _06107_ | _06106_;
  assign _06109_ = sel_oi_one_hot_i[210] & i[33];
  assign _06110_ = sel_oi_one_hot_i[211] & i[49];
  assign _06111_ = _06110_ | _06109_;
  assign _06112_ = _06111_ | _06108_;
  assign _06113_ = sel_oi_one_hot_i[212] & i[65];
  assign _06114_ = sel_oi_one_hot_i[213] & i[81];
  assign _06115_ = _06114_ | _06113_;
  assign _06116_ = sel_oi_one_hot_i[214] & i[97];
  assign _06117_ = sel_oi_one_hot_i[215] & i[113];
  assign _06118_ = _06117_ | _06116_;
  assign _06119_ = _06118_ | _06115_;
  assign _06120_ = _06119_ | _06112_;
  assign _06121_ = sel_oi_one_hot_i[216] & i[129];
  assign _06122_ = sel_oi_one_hot_i[217] & i[145];
  assign _06123_ = _06122_ | _06121_;
  assign _06124_ = sel_oi_one_hot_i[218] & i[161];
  assign _06125_ = sel_oi_one_hot_i[219] & i[177];
  assign _06126_ = _06125_ | _06124_;
  assign _06127_ = _06126_ | _06123_;
  assign _06128_ = sel_oi_one_hot_i[220] & i[193];
  assign _06129_ = sel_oi_one_hot_i[221] & i[209];
  assign _06130_ = _06129_ | _06128_;
  assign _06131_ = sel_oi_one_hot_i[222] & i[225];
  assign _06132_ = sel_oi_one_hot_i[223] & i[241];
  assign _06133_ = _06132_ | _06131_;
  assign _06134_ = _06133_ | _06130_;
  assign _06135_ = _06134_ | _06127_;
  assign o[209] = _06135_ | _06120_;
  assign _06136_ = sel_oi_one_hot_i[208] & i[0];
  assign _06137_ = sel_oi_one_hot_i[209] & i[16];
  assign _06138_ = _06137_ | _06136_;
  assign _06139_ = sel_oi_one_hot_i[210] & i[32];
  assign _06140_ = sel_oi_one_hot_i[211] & i[48];
  assign _06141_ = _06140_ | _06139_;
  assign _06142_ = _06141_ | _06138_;
  assign _06143_ = sel_oi_one_hot_i[212] & i[64];
  assign _06144_ = sel_oi_one_hot_i[213] & i[80];
  assign _06145_ = _06144_ | _06143_;
  assign _06146_ = sel_oi_one_hot_i[214] & i[96];
  assign _06147_ = sel_oi_one_hot_i[215] & i[112];
  assign _06148_ = _06147_ | _06146_;
  assign _06149_ = _06148_ | _06145_;
  assign _06150_ = _06149_ | _06142_;
  assign _06151_ = sel_oi_one_hot_i[216] & i[128];
  assign _06152_ = sel_oi_one_hot_i[217] & i[144];
  assign _06153_ = _06152_ | _06151_;
  assign _06154_ = sel_oi_one_hot_i[218] & i[160];
  assign _06155_ = sel_oi_one_hot_i[219] & i[176];
  assign _06156_ = _06155_ | _06154_;
  assign _06157_ = _06156_ | _06153_;
  assign _06158_ = sel_oi_one_hot_i[220] & i[192];
  assign _06159_ = sel_oi_one_hot_i[221] & i[208];
  assign _06160_ = _06159_ | _06158_;
  assign _06161_ = sel_oi_one_hot_i[222] & i[224];
  assign _06162_ = sel_oi_one_hot_i[223] & i[240];
  assign _06163_ = _06162_ | _06161_;
  assign _06164_ = _06163_ | _06160_;
  assign _06165_ = _06164_ | _06157_;
  assign o[208] = _06165_ | _06150_;
  assign _06166_ = i[10] & sel_oi_one_hot_i[16];
  assign _06167_ = i[26] & sel_oi_one_hot_i[17];
  assign _06168_ = _06167_ | _06166_;
  assign _06169_ = i[42] & sel_oi_one_hot_i[18];
  assign _06170_ = i[58] & sel_oi_one_hot_i[19];
  assign _06171_ = _06170_ | _06169_;
  assign _06172_ = _06171_ | _06168_;
  assign _06173_ = i[74] & sel_oi_one_hot_i[20];
  assign _06174_ = i[90] & sel_oi_one_hot_i[21];
  assign _06175_ = _06174_ | _06173_;
  assign _06176_ = i[106] & sel_oi_one_hot_i[22];
  assign _06177_ = i[122] & sel_oi_one_hot_i[23];
  assign _06178_ = _06177_ | _06176_;
  assign _06179_ = _06178_ | _06175_;
  assign _06180_ = _06179_ | _06172_;
  assign _06181_ = i[138] & sel_oi_one_hot_i[24];
  assign _06182_ = i[154] & sel_oi_one_hot_i[25];
  assign _06183_ = _06182_ | _06181_;
  assign _06184_ = i[170] & sel_oi_one_hot_i[26];
  assign _06185_ = i[186] & sel_oi_one_hot_i[27];
  assign _06186_ = _06185_ | _06184_;
  assign _06187_ = _06186_ | _06183_;
  assign _06188_ = i[202] & sel_oi_one_hot_i[28];
  assign _06189_ = i[218] & sel_oi_one_hot_i[29];
  assign _06190_ = _06189_ | _06188_;
  assign _06191_ = sel_oi_one_hot_i[30] & i[234];
  assign _06192_ = sel_oi_one_hot_i[31] & i[250];
  assign _06193_ = _06192_ | _06191_;
  assign _06194_ = _06193_ | _06190_;
  assign _06195_ = _06194_ | _06187_;
  assign o[26] = _06195_ | _06180_;
  assign _06196_ = sel_oi_one_hot_i[224] & i[15];
  assign _06197_ = sel_oi_one_hot_i[225] & i[31];
  assign _06198_ = _06197_ | _06196_;
  assign _06199_ = sel_oi_one_hot_i[226] & i[47];
  assign _06200_ = sel_oi_one_hot_i[227] & i[63];
  assign _06201_ = _06200_ | _06199_;
  assign _06202_ = _06201_ | _06198_;
  assign _06203_ = sel_oi_one_hot_i[228] & i[79];
  assign _06204_ = sel_oi_one_hot_i[229] & i[95];
  assign _06205_ = _06204_ | _06203_;
  assign _06206_ = sel_oi_one_hot_i[230] & i[111];
  assign _06207_ = sel_oi_one_hot_i[231] & i[127];
  assign _06208_ = _06207_ | _06206_;
  assign _06209_ = _06208_ | _06205_;
  assign _06210_ = _06209_ | _06202_;
  assign _06211_ = sel_oi_one_hot_i[232] & i[143];
  assign _06212_ = sel_oi_one_hot_i[233] & i[159];
  assign _06213_ = _06212_ | _06211_;
  assign _06214_ = sel_oi_one_hot_i[234] & i[175];
  assign _06215_ = sel_oi_one_hot_i[235] & i[191];
  assign _06216_ = _06215_ | _06214_;
  assign _06217_ = _06216_ | _06213_;
  assign _06218_ = sel_oi_one_hot_i[236] & i[207];
  assign _06219_ = sel_oi_one_hot_i[237] & i[223];
  assign _06220_ = _06219_ | _06218_;
  assign _06221_ = sel_oi_one_hot_i[238] & i[239];
  assign _06222_ = sel_oi_one_hot_i[239] & i[255];
  assign _06223_ = _06222_ | _06221_;
  assign _06224_ = _06223_ | _06220_;
  assign _06225_ = _06224_ | _06217_;
  assign o[239] = _06225_ | _06210_;
  assign _06226_ = sel_oi_one_hot_i[224] & i[14];
  assign _06227_ = sel_oi_one_hot_i[225] & i[30];
  assign _06228_ = _06227_ | _06226_;
  assign _06229_ = sel_oi_one_hot_i[226] & i[46];
  assign _06230_ = sel_oi_one_hot_i[227] & i[62];
  assign _06231_ = _06230_ | _06229_;
  assign _06232_ = _06231_ | _06228_;
  assign _06233_ = sel_oi_one_hot_i[228] & i[78];
  assign _06234_ = sel_oi_one_hot_i[229] & i[94];
  assign _06235_ = _06234_ | _06233_;
  assign _06236_ = sel_oi_one_hot_i[230] & i[110];
  assign _06237_ = sel_oi_one_hot_i[231] & i[126];
  assign _06238_ = _06237_ | _06236_;
  assign _06239_ = _06238_ | _06235_;
  assign _06240_ = _06239_ | _06232_;
  assign _06241_ = sel_oi_one_hot_i[232] & i[142];
  assign _06242_ = sel_oi_one_hot_i[233] & i[158];
  assign _06243_ = _06242_ | _06241_;
  assign _06244_ = sel_oi_one_hot_i[234] & i[174];
  assign _06245_ = sel_oi_one_hot_i[235] & i[190];
  assign _06246_ = _06245_ | _06244_;
  assign _06247_ = _06246_ | _06243_;
  assign _06248_ = sel_oi_one_hot_i[236] & i[206];
  assign _06249_ = sel_oi_one_hot_i[237] & i[222];
  assign _06250_ = _06249_ | _06248_;
  assign _06251_ = sel_oi_one_hot_i[238] & i[238];
  assign _06252_ = sel_oi_one_hot_i[239] & i[254];
  assign _06253_ = _06252_ | _06251_;
  assign _06254_ = _06253_ | _06250_;
  assign _06255_ = _06254_ | _06247_;
  assign o[238] = _06255_ | _06240_;
  assign _06256_ = sel_oi_one_hot_i[224] & i[13];
  assign _06257_ = sel_oi_one_hot_i[225] & i[29];
  assign _06258_ = _06257_ | _06256_;
  assign _06259_ = sel_oi_one_hot_i[226] & i[45];
  assign _06260_ = sel_oi_one_hot_i[227] & i[61];
  assign _06261_ = _06260_ | _06259_;
  assign _06262_ = _06261_ | _06258_;
  assign _06263_ = sel_oi_one_hot_i[228] & i[77];
  assign _06264_ = sel_oi_one_hot_i[229] & i[93];
  assign _06265_ = _06264_ | _06263_;
  assign _06266_ = sel_oi_one_hot_i[230] & i[109];
  assign _06267_ = sel_oi_one_hot_i[231] & i[125];
  assign _06268_ = _06267_ | _06266_;
  assign _06269_ = _06268_ | _06265_;
  assign _06270_ = _06269_ | _06262_;
  assign _06271_ = sel_oi_one_hot_i[232] & i[141];
  assign _06272_ = sel_oi_one_hot_i[233] & i[157];
  assign _06273_ = _06272_ | _06271_;
  assign _06274_ = sel_oi_one_hot_i[234] & i[173];
  assign _06275_ = sel_oi_one_hot_i[235] & i[189];
  assign _06276_ = _06275_ | _06274_;
  assign _06277_ = _06276_ | _06273_;
  assign _06278_ = sel_oi_one_hot_i[236] & i[205];
  assign _06279_ = sel_oi_one_hot_i[237] & i[221];
  assign _06280_ = _06279_ | _06278_;
  assign _06281_ = sel_oi_one_hot_i[238] & i[237];
  assign _06282_ = sel_oi_one_hot_i[239] & i[253];
  assign _06283_ = _06282_ | _06281_;
  assign _06284_ = _06283_ | _06280_;
  assign _06285_ = _06284_ | _06277_;
  assign o[237] = _06285_ | _06270_;
  assign _06286_ = i[9] & sel_oi_one_hot_i[16];
  assign _06287_ = i[25] & sel_oi_one_hot_i[17];
  assign _06288_ = _06287_ | _06286_;
  assign _06289_ = i[41] & sel_oi_one_hot_i[18];
  assign _06290_ = i[57] & sel_oi_one_hot_i[19];
  assign _06291_ = _06290_ | _06289_;
  assign _06292_ = _06291_ | _06288_;
  assign _06293_ = i[73] & sel_oi_one_hot_i[20];
  assign _06294_ = i[89] & sel_oi_one_hot_i[21];
  assign _06295_ = _06294_ | _06293_;
  assign _06296_ = i[105] & sel_oi_one_hot_i[22];
  assign _06297_ = i[121] & sel_oi_one_hot_i[23];
  assign _06298_ = _06297_ | _06296_;
  assign _06299_ = _06298_ | _06295_;
  assign _06300_ = _06299_ | _06292_;
  assign _06301_ = i[137] & sel_oi_one_hot_i[24];
  assign _06302_ = i[153] & sel_oi_one_hot_i[25];
  assign _06303_ = _06302_ | _06301_;
  assign _06304_ = i[169] & sel_oi_one_hot_i[26];
  assign _06305_ = i[185] & sel_oi_one_hot_i[27];
  assign _06306_ = _06305_ | _06304_;
  assign _06307_ = _06306_ | _06303_;
  assign _06308_ = i[201] & sel_oi_one_hot_i[28];
  assign _06309_ = i[217] & sel_oi_one_hot_i[29];
  assign _06310_ = _06309_ | _06308_;
  assign _06311_ = i[233] & sel_oi_one_hot_i[30];
  assign _06312_ = sel_oi_one_hot_i[31] & i[249];
  assign _06313_ = _06312_ | _06311_;
  assign _06314_ = _06313_ | _06310_;
  assign _06315_ = _06314_ | _06307_;
  assign o[25] = _06315_ | _06300_;
  assign _06316_ = sel_oi_one_hot_i[224] & i[12];
  assign _06317_ = sel_oi_one_hot_i[225] & i[28];
  assign _06318_ = _06317_ | _06316_;
  assign _06319_ = sel_oi_one_hot_i[226] & i[44];
  assign _06320_ = sel_oi_one_hot_i[227] & i[60];
  assign _06321_ = _06320_ | _06319_;
  assign _06322_ = _06321_ | _06318_;
  assign _06323_ = sel_oi_one_hot_i[228] & i[76];
  assign _06324_ = sel_oi_one_hot_i[229] & i[92];
  assign _06325_ = _06324_ | _06323_;
  assign _06326_ = sel_oi_one_hot_i[230] & i[108];
  assign _06327_ = sel_oi_one_hot_i[231] & i[124];
  assign _06328_ = _06327_ | _06326_;
  assign _06329_ = _06328_ | _06325_;
  assign _06330_ = _06329_ | _06322_;
  assign _06331_ = sel_oi_one_hot_i[232] & i[140];
  assign _06332_ = sel_oi_one_hot_i[233] & i[156];
  assign _06333_ = _06332_ | _06331_;
  assign _06334_ = sel_oi_one_hot_i[234] & i[172];
  assign _06335_ = sel_oi_one_hot_i[235] & i[188];
  assign _06336_ = _06335_ | _06334_;
  assign _06337_ = _06336_ | _06333_;
  assign _06338_ = sel_oi_one_hot_i[236] & i[204];
  assign _06339_ = sel_oi_one_hot_i[237] & i[220];
  assign _06340_ = _06339_ | _06338_;
  assign _06341_ = sel_oi_one_hot_i[238] & i[236];
  assign _06342_ = sel_oi_one_hot_i[239] & i[252];
  assign _06343_ = _06342_ | _06341_;
  assign _06344_ = _06343_ | _06340_;
  assign _06345_ = _06344_ | _06337_;
  assign o[236] = _06345_ | _06330_;
  assign _06346_ = sel_oi_one_hot_i[224] & i[11];
  assign _06347_ = sel_oi_one_hot_i[225] & i[27];
  assign _06348_ = _06347_ | _06346_;
  assign _06349_ = sel_oi_one_hot_i[226] & i[43];
  assign _06350_ = sel_oi_one_hot_i[227] & i[59];
  assign _06351_ = _06350_ | _06349_;
  assign _06352_ = _06351_ | _06348_;
  assign _06353_ = sel_oi_one_hot_i[228] & i[75];
  assign _06354_ = sel_oi_one_hot_i[229] & i[91];
  assign _06355_ = _06354_ | _06353_;
  assign _06356_ = sel_oi_one_hot_i[230] & i[107];
  assign _06357_ = sel_oi_one_hot_i[231] & i[123];
  assign _06358_ = _06357_ | _06356_;
  assign _06359_ = _06358_ | _06355_;
  assign _06360_ = _06359_ | _06352_;
  assign _06361_ = sel_oi_one_hot_i[232] & i[139];
  assign _06362_ = sel_oi_one_hot_i[233] & i[155];
  assign _06363_ = _06362_ | _06361_;
  assign _06364_ = sel_oi_one_hot_i[234] & i[171];
  assign _06365_ = sel_oi_one_hot_i[235] & i[187];
  assign _06366_ = _06365_ | _06364_;
  assign _06367_ = _06366_ | _06363_;
  assign _06368_ = sel_oi_one_hot_i[236] & i[203];
  assign _06369_ = sel_oi_one_hot_i[237] & i[219];
  assign _06370_ = _06369_ | _06368_;
  assign _06371_ = sel_oi_one_hot_i[238] & i[235];
  assign _06372_ = sel_oi_one_hot_i[239] & i[251];
  assign _06373_ = _06372_ | _06371_;
  assign _06374_ = _06373_ | _06370_;
  assign _06375_ = _06374_ | _06367_;
  assign o[235] = _06375_ | _06360_;
  assign _06376_ = sel_oi_one_hot_i[224] & i[10];
  assign _06377_ = sel_oi_one_hot_i[225] & i[26];
  assign _06378_ = _06377_ | _06376_;
  assign _06379_ = sel_oi_one_hot_i[226] & i[42];
  assign _06380_ = sel_oi_one_hot_i[227] & i[58];
  assign _06381_ = _06380_ | _06379_;
  assign _06382_ = _06381_ | _06378_;
  assign _06383_ = sel_oi_one_hot_i[228] & i[74];
  assign _06384_ = sel_oi_one_hot_i[229] & i[90];
  assign _06385_ = _06384_ | _06383_;
  assign _06386_ = sel_oi_one_hot_i[230] & i[106];
  assign _06387_ = sel_oi_one_hot_i[231] & i[122];
  assign _06388_ = _06387_ | _06386_;
  assign _06389_ = _06388_ | _06385_;
  assign _06390_ = _06389_ | _06382_;
  assign _06391_ = sel_oi_one_hot_i[232] & i[138];
  assign _06392_ = sel_oi_one_hot_i[233] & i[154];
  assign _06393_ = _06392_ | _06391_;
  assign _06394_ = sel_oi_one_hot_i[234] & i[170];
  assign _06395_ = sel_oi_one_hot_i[235] & i[186];
  assign _06396_ = _06395_ | _06394_;
  assign _06397_ = _06396_ | _06393_;
  assign _06398_ = sel_oi_one_hot_i[236] & i[202];
  assign _06399_ = sel_oi_one_hot_i[237] & i[218];
  assign _06400_ = _06399_ | _06398_;
  assign _06401_ = sel_oi_one_hot_i[238] & i[234];
  assign _06402_ = sel_oi_one_hot_i[239] & i[250];
  assign _06403_ = _06402_ | _06401_;
  assign _06404_ = _06403_ | _06400_;
  assign _06405_ = _06404_ | _06397_;
  assign o[234] = _06405_ | _06390_;
  assign _06406_ = sel_oi_one_hot_i[224] & i[9];
  assign _06407_ = sel_oi_one_hot_i[225] & i[25];
  assign _06408_ = _06407_ | _06406_;
  assign _06409_ = sel_oi_one_hot_i[226] & i[41];
  assign _06410_ = sel_oi_one_hot_i[227] & i[57];
  assign _06411_ = _06410_ | _06409_;
  assign _06412_ = _06411_ | _06408_;
  assign _06413_ = sel_oi_one_hot_i[228] & i[73];
  assign _06414_ = sel_oi_one_hot_i[229] & i[89];
  assign _06415_ = _06414_ | _06413_;
  assign _06416_ = sel_oi_one_hot_i[230] & i[105];
  assign _06417_ = sel_oi_one_hot_i[231] & i[121];
  assign _06418_ = _06417_ | _06416_;
  assign _06419_ = _06418_ | _06415_;
  assign _06420_ = _06419_ | _06412_;
  assign _06421_ = sel_oi_one_hot_i[232] & i[137];
  assign _06422_ = sel_oi_one_hot_i[233] & i[153];
  assign _06423_ = _06422_ | _06421_;
  assign _06424_ = sel_oi_one_hot_i[234] & i[169];
  assign _06425_ = sel_oi_one_hot_i[235] & i[185];
  assign _06426_ = _06425_ | _06424_;
  assign _06427_ = _06426_ | _06423_;
  assign _06428_ = sel_oi_one_hot_i[236] & i[201];
  assign _06429_ = sel_oi_one_hot_i[237] & i[217];
  assign _06430_ = _06429_ | _06428_;
  assign _06431_ = sel_oi_one_hot_i[238] & i[233];
  assign _06432_ = sel_oi_one_hot_i[239] & i[249];
  assign _06433_ = _06432_ | _06431_;
  assign _06434_ = _06433_ | _06430_;
  assign _06435_ = _06434_ | _06427_;
  assign o[233] = _06435_ | _06420_;
  assign _06436_ = sel_oi_one_hot_i[224] & i[8];
  assign _06437_ = sel_oi_one_hot_i[225] & i[24];
  assign _06438_ = _06437_ | _06436_;
  assign _06439_ = sel_oi_one_hot_i[226] & i[40];
  assign _06440_ = sel_oi_one_hot_i[227] & i[56];
  assign _06441_ = _06440_ | _06439_;
  assign _06442_ = _06441_ | _06438_;
  assign _06443_ = sel_oi_one_hot_i[228] & i[72];
  assign _06444_ = sel_oi_one_hot_i[229] & i[88];
  assign _06445_ = _06444_ | _06443_;
  assign _06446_ = sel_oi_one_hot_i[230] & i[104];
  assign _06447_ = sel_oi_one_hot_i[231] & i[120];
  assign _06448_ = _06447_ | _06446_;
  assign _06449_ = _06448_ | _06445_;
  assign _06450_ = _06449_ | _06442_;
  assign _06451_ = sel_oi_one_hot_i[232] & i[136];
  assign _06452_ = sel_oi_one_hot_i[233] & i[152];
  assign _06453_ = _06452_ | _06451_;
  assign _06454_ = sel_oi_one_hot_i[234] & i[168];
  assign _06455_ = sel_oi_one_hot_i[235] & i[184];
  assign _06456_ = _06455_ | _06454_;
  assign _06457_ = _06456_ | _06453_;
  assign _06458_ = sel_oi_one_hot_i[236] & i[200];
  assign _06459_ = sel_oi_one_hot_i[237] & i[216];
  assign _06460_ = _06459_ | _06458_;
  assign _06461_ = sel_oi_one_hot_i[238] & i[232];
  assign _06462_ = sel_oi_one_hot_i[239] & i[248];
  assign _06463_ = _06462_ | _06461_;
  assign _06464_ = _06463_ | _06460_;
  assign _06465_ = _06464_ | _06457_;
  assign o[232] = _06465_ | _06450_;
  assign _06466_ = sel_oi_one_hot_i[224] & i[7];
  assign _06467_ = sel_oi_one_hot_i[225] & i[23];
  assign _06468_ = _06467_ | _06466_;
  assign _06469_ = sel_oi_one_hot_i[226] & i[39];
  assign _06470_ = sel_oi_one_hot_i[227] & i[55];
  assign _06471_ = _06470_ | _06469_;
  assign _06472_ = _06471_ | _06468_;
  assign _06473_ = sel_oi_one_hot_i[228] & i[71];
  assign _06474_ = sel_oi_one_hot_i[229] & i[87];
  assign _06475_ = _06474_ | _06473_;
  assign _06476_ = sel_oi_one_hot_i[230] & i[103];
  assign _06477_ = sel_oi_one_hot_i[231] & i[119];
  assign _06478_ = _06477_ | _06476_;
  assign _06479_ = _06478_ | _06475_;
  assign _06480_ = _06479_ | _06472_;
  assign _06481_ = sel_oi_one_hot_i[232] & i[135];
  assign _06482_ = sel_oi_one_hot_i[233] & i[151];
  assign _06483_ = _06482_ | _06481_;
  assign _06485_ = sel_oi_one_hot_i[234] & i[167];
  assign _06486_ = sel_oi_one_hot_i[235] & i[183];
  assign _06487_ = _06486_ | _06485_;
  assign _06488_ = _06487_ | _06483_;
  assign _06489_ = sel_oi_one_hot_i[236] & i[199];
  assign _06490_ = sel_oi_one_hot_i[237] & i[215];
  assign _06491_ = _06490_ | _06489_;
  assign _06492_ = sel_oi_one_hot_i[238] & i[231];
  assign _06493_ = sel_oi_one_hot_i[239] & i[247];
  assign _06494_ = _06493_ | _06492_;
  assign _06496_ = _06494_ | _06491_;
  assign _06497_ = _06496_ | _06488_;
  assign o[231] = _06497_ | _06480_;
  assign _06498_ = sel_oi_one_hot_i[224] & i[6];
  assign _06499_ = sel_oi_one_hot_i[225] & i[22];
  assign _06500_ = _06499_ | _06498_;
  assign _06501_ = sel_oi_one_hot_i[226] & i[38];
  assign _06502_ = sel_oi_one_hot_i[227] & i[54];
  assign _06503_ = _06502_ | _06501_;
  assign _06504_ = _06503_ | _06500_;
  assign _06506_ = sel_oi_one_hot_i[228] & i[70];
  assign _06507_ = sel_oi_one_hot_i[229] & i[86];
  assign _06508_ = _06507_ | _06506_;
  assign _06509_ = sel_oi_one_hot_i[230] & i[102];
  assign _06510_ = sel_oi_one_hot_i[231] & i[118];
  assign _06511_ = _06510_ | _06509_;
  assign _06512_ = _06511_ | _06508_;
  assign _06513_ = _06512_ | _06504_;
  assign _06514_ = sel_oi_one_hot_i[232] & i[134];
  assign _06515_ = sel_oi_one_hot_i[233] & i[150];
  assign _06517_ = _06515_ | _06514_;
  assign _06518_ = sel_oi_one_hot_i[234] & i[166];
  assign _06519_ = sel_oi_one_hot_i[235] & i[182];
  assign _06520_ = _06519_ | _06518_;
  assign _06521_ = _06520_ | _06517_;
  assign _06522_ = sel_oi_one_hot_i[236] & i[198];
  assign _06523_ = sel_oi_one_hot_i[237] & i[214];
  assign _06524_ = _06523_ | _06522_;
  assign _06525_ = sel_oi_one_hot_i[238] & i[230];
  assign _06526_ = sel_oi_one_hot_i[239] & i[246];
  assign _06528_ = _06526_ | _06525_;
  assign _06529_ = _06528_ | _06524_;
  assign _06530_ = _06529_ | _06521_;
  assign o[230] = _06530_ | _06513_;
  assign _06531_ = sel_oi_one_hot_i[224] & i[5];
  assign _06532_ = sel_oi_one_hot_i[225] & i[21];
  assign _06533_ = _06532_ | _06531_;
  assign _06534_ = sel_oi_one_hot_i[226] & i[37];
  assign _06535_ = sel_oi_one_hot_i[227] & i[53];
  assign _06536_ = _06535_ | _06534_;
  assign _06538_ = _06536_ | _06533_;
  assign _06539_ = sel_oi_one_hot_i[228] & i[69];
  assign _06540_ = sel_oi_one_hot_i[229] & i[85];
  assign _06541_ = _06540_ | _06539_;
  assign _06542_ = sel_oi_one_hot_i[230] & i[101];
  assign _06543_ = sel_oi_one_hot_i[231] & i[117];
  assign _06544_ = _06543_ | _06542_;
  assign _06545_ = _06544_ | _06541_;
  assign _06546_ = _06545_ | _06538_;
  assign _06547_ = sel_oi_one_hot_i[232] & i[133];
  assign _06549_ = sel_oi_one_hot_i[233] & i[149];
  assign _06550_ = _06549_ | _06547_;
  assign _06551_ = sel_oi_one_hot_i[234] & i[165];
  assign _06552_ = sel_oi_one_hot_i[235] & i[181];
  assign _06553_ = _06552_ | _06551_;
  assign _06554_ = _06553_ | _06550_;
  assign _06555_ = sel_oi_one_hot_i[236] & i[197];
  assign _06556_ = sel_oi_one_hot_i[237] & i[213];
  assign _06557_ = _06556_ | _06555_;
  assign _06558_ = sel_oi_one_hot_i[238] & i[229];
  assign _06560_ = sel_oi_one_hot_i[239] & i[245];
  assign _06561_ = _06560_ | _06558_;
  assign _06562_ = _06561_ | _06557_;
  assign _06563_ = _06562_ | _06554_;
  assign o[229] = _06563_ | _06546_;
  assign _06564_ = sel_oi_one_hot_i[224] & i[4];
  assign _06565_ = sel_oi_one_hot_i[225] & i[20];
  assign _06566_ = _06565_ | _06564_;
  assign _06567_ = sel_oi_one_hot_i[226] & i[36];
  assign _06568_ = sel_oi_one_hot_i[227] & i[52];
  assign _06570_ = _06568_ | _06567_;
  assign _06571_ = _06570_ | _06566_;
  assign _06572_ = sel_oi_one_hot_i[228] & i[68];
  assign _06573_ = sel_oi_one_hot_i[229] & i[84];
  assign _06574_ = _06573_ | _06572_;
  assign _06575_ = sel_oi_one_hot_i[230] & i[100];
  assign _06576_ = sel_oi_one_hot_i[231] & i[116];
  assign _06577_ = _06576_ | _06575_;
  assign _06578_ = _06577_ | _06574_;
  assign _06579_ = _06578_ | _06571_;
  assign _06581_ = sel_oi_one_hot_i[232] & i[132];
  assign _06582_ = sel_oi_one_hot_i[233] & i[148];
  assign _06583_ = _06582_ | _06581_;
  assign _06584_ = sel_oi_one_hot_i[234] & i[164];
  assign _06585_ = sel_oi_one_hot_i[235] & i[180];
  assign _06586_ = _06585_ | _06584_;
  assign _06587_ = _06586_ | _06583_;
  assign _06588_ = sel_oi_one_hot_i[236] & i[196];
  assign _06589_ = sel_oi_one_hot_i[237] & i[212];
  assign _06590_ = _06589_ | _06588_;
  assign _06592_ = sel_oi_one_hot_i[238] & i[228];
  assign _06593_ = sel_oi_one_hot_i[239] & i[244];
  assign _06594_ = _06593_ | _06592_;
  assign _06595_ = _06594_ | _06590_;
  assign _06596_ = _06595_ | _06587_;
  assign o[228] = _06596_ | _06579_;
  assign _06597_ = sel_oi_one_hot_i[224] & i[3];
  assign _06598_ = sel_oi_one_hot_i[225] & i[19];
  assign _06599_ = _06598_ | _06597_;
  assign _06600_ = sel_oi_one_hot_i[226] & i[35];
  assign _06602_ = sel_oi_one_hot_i[227] & i[51];
  assign _06603_ = _06602_ | _06600_;
  assign _06604_ = _06603_ | _06599_;
  assign _06605_ = sel_oi_one_hot_i[228] & i[67];
  assign _06606_ = sel_oi_one_hot_i[229] & i[83];
  assign _06607_ = _06606_ | _06605_;
  assign _06608_ = sel_oi_one_hot_i[230] & i[99];
  assign _06609_ = sel_oi_one_hot_i[231] & i[115];
  assign _06610_ = _06609_ | _06608_;
  assign _06611_ = _06610_ | _06607_;
  assign _06613_ = _06611_ | _06604_;
  assign _06614_ = sel_oi_one_hot_i[232] & i[131];
  assign _06615_ = sel_oi_one_hot_i[233] & i[147];
  assign _06616_ = _06615_ | _06614_;
  assign _06617_ = sel_oi_one_hot_i[234] & i[163];
  assign _06618_ = sel_oi_one_hot_i[235] & i[179];
  assign _06619_ = _06618_ | _06617_;
  assign _06620_ = _06619_ | _06616_;
  assign _06621_ = sel_oi_one_hot_i[236] & i[195];
  assign _06622_ = sel_oi_one_hot_i[237] & i[211];
  assign _06624_ = _06622_ | _06621_;
  assign _06625_ = sel_oi_one_hot_i[238] & i[227];
  assign _06626_ = sel_oi_one_hot_i[239] & i[243];
  assign _06627_ = _06626_ | _06625_;
  assign _06628_ = _06627_ | _06624_;
  assign _06629_ = _06628_ | _06620_;
  assign o[227] = _06629_ | _06613_;
  assign _06630_ = i[8] & sel_oi_one_hot_i[16];
  assign _06631_ = i[24] & sel_oi_one_hot_i[17];
  assign _06632_ = _06631_ | _06630_;
  assign _06634_ = i[40] & sel_oi_one_hot_i[18];
  assign _06635_ = i[56] & sel_oi_one_hot_i[19];
  assign _06636_ = _06635_ | _06634_;
  assign _06637_ = _06636_ | _06632_;
  assign _06638_ = i[72] & sel_oi_one_hot_i[20];
  assign _06639_ = i[88] & sel_oi_one_hot_i[21];
  assign _06640_ = _06639_ | _06638_;
  assign _06641_ = i[104] & sel_oi_one_hot_i[22];
  assign _06642_ = i[120] & sel_oi_one_hot_i[23];
  assign _06643_ = _06642_ | _06641_;
  assign _06645_ = _06643_ | _06640_;
  assign _06646_ = _06645_ | _06637_;
  assign _06647_ = i[136] & sel_oi_one_hot_i[24];
  assign _06648_ = i[152] & sel_oi_one_hot_i[25];
  assign _06649_ = _06648_ | _06647_;
  assign _06650_ = i[168] & sel_oi_one_hot_i[26];
  assign _06651_ = i[184] & sel_oi_one_hot_i[27];
  assign _06652_ = _06651_ | _06650_;
  assign _06653_ = _06652_ | _06649_;
  assign _06654_ = i[200] & sel_oi_one_hot_i[28];
  assign _06656_ = i[216] & sel_oi_one_hot_i[29];
  assign _06657_ = _06656_ | _06654_;
  assign _06658_ = i[232] & sel_oi_one_hot_i[30];
  assign _06659_ = sel_oi_one_hot_i[31] & i[248];
  assign _06660_ = _06659_ | _06658_;
  assign _06661_ = _06660_ | _06657_;
  assign _06662_ = _06661_ | _06653_;
  assign o[24] = _06662_ | _06646_;
  assign _06663_ = sel_oi_one_hot_i[224] & i[2];
  assign _06664_ = sel_oi_one_hot_i[225] & i[18];
  assign _06666_ = _06664_ | _06663_;
  assign _06667_ = sel_oi_one_hot_i[226] & i[34];
  assign _06668_ = sel_oi_one_hot_i[227] & i[50];
  assign _06669_ = _06668_ | _06667_;
  assign _06670_ = _06669_ | _06666_;
  assign _06671_ = sel_oi_one_hot_i[228] & i[66];
  assign _06672_ = sel_oi_one_hot_i[229] & i[82];
  assign _06673_ = _06672_ | _06671_;
  assign _06674_ = sel_oi_one_hot_i[230] & i[98];
  assign _06675_ = sel_oi_one_hot_i[231] & i[114];
  assign _06677_ = _06675_ | _06674_;
  assign _06678_ = _06677_ | _06673_;
  assign _06679_ = _06678_ | _06670_;
  assign _06680_ = sel_oi_one_hot_i[232] & i[130];
  assign _06681_ = sel_oi_one_hot_i[233] & i[146];
  assign _06682_ = _06681_ | _06680_;
  assign _06683_ = sel_oi_one_hot_i[234] & i[162];
  assign _06684_ = sel_oi_one_hot_i[235] & i[178];
  assign _06685_ = _06684_ | _06683_;
  assign _06686_ = _06685_ | _06682_;
  assign _06688_ = sel_oi_one_hot_i[236] & i[194];
  assign _06689_ = sel_oi_one_hot_i[237] & i[210];
  assign _06690_ = _06689_ | _06688_;
  assign _06691_ = sel_oi_one_hot_i[238] & i[226];
  assign _06692_ = sel_oi_one_hot_i[239] & i[242];
  assign _06693_ = _06692_ | _06691_;
  assign _06694_ = _06693_ | _06690_;
  assign _06695_ = _06694_ | _06686_;
  assign o[226] = _06695_ | _06679_;
  assign _06696_ = sel_oi_one_hot_i[224] & i[1];
  assign _06698_ = sel_oi_one_hot_i[225] & i[17];
  assign _06699_ = _06698_ | _06696_;
  assign _06700_ = sel_oi_one_hot_i[226] & i[33];
  assign _06701_ = sel_oi_one_hot_i[227] & i[49];
  assign _06702_ = _06701_ | _06700_;
  assign _06703_ = _06702_ | _06699_;
  assign _06704_ = sel_oi_one_hot_i[228] & i[65];
  assign _06705_ = sel_oi_one_hot_i[229] & i[81];
  assign _06706_ = _06705_ | _06704_;
  assign _06707_ = sel_oi_one_hot_i[230] & i[97];
  assign _06709_ = sel_oi_one_hot_i[231] & i[113];
  assign _06710_ = _06709_ | _06707_;
  assign _06711_ = _06710_ | _06706_;
  assign _06712_ = _06711_ | _06703_;
  assign _06713_ = sel_oi_one_hot_i[232] & i[129];
  assign _06714_ = sel_oi_one_hot_i[233] & i[145];
  assign _06715_ = _06714_ | _06713_;
  assign _06716_ = sel_oi_one_hot_i[234] & i[161];
  assign _06717_ = sel_oi_one_hot_i[235] & i[177];
  assign _06718_ = _06717_ | _06716_;
  assign _06720_ = _06718_ | _06715_;
  assign _06721_ = sel_oi_one_hot_i[236] & i[193];
  assign _06722_ = sel_oi_one_hot_i[237] & i[209];
  assign _06723_ = _06722_ | _06721_;
  assign _06724_ = sel_oi_one_hot_i[238] & i[225];
  assign _06725_ = sel_oi_one_hot_i[239] & i[241];
  assign _06726_ = _06725_ | _06724_;
  assign _06727_ = _06726_ | _06723_;
  assign _06728_ = _06727_ | _06720_;
  assign o[225] = _06728_ | _06712_;
  assign _06730_ = sel_oi_one_hot_i[224] & i[0];
  assign _06731_ = sel_oi_one_hot_i[225] & i[16];
  assign _06732_ = _06731_ | _06730_;
  assign _06733_ = sel_oi_one_hot_i[226] & i[32];
  assign _06734_ = sel_oi_one_hot_i[227] & i[48];
  assign _06735_ = _06734_ | _06733_;
  assign _06736_ = _06735_ | _06732_;
  assign _06737_ = sel_oi_one_hot_i[228] & i[64];
  assign _06738_ = sel_oi_one_hot_i[229] & i[80];
  assign _06739_ = _06738_ | _06737_;
  assign _06741_ = sel_oi_one_hot_i[230] & i[96];
  assign _06742_ = sel_oi_one_hot_i[231] & i[112];
  assign _06743_ = _06742_ | _06741_;
  assign _06744_ = _06743_ | _06739_;
  assign _06745_ = _06744_ | _06736_;
  assign _06746_ = sel_oi_one_hot_i[232] & i[128];
  assign _06747_ = sel_oi_one_hot_i[233] & i[144];
  assign _06748_ = _06747_ | _06746_;
  assign _06749_ = sel_oi_one_hot_i[234] & i[160];
  assign _06750_ = sel_oi_one_hot_i[235] & i[176];
  assign _06752_ = _06750_ | _06749_;
  assign _06753_ = _06752_ | _06748_;
  assign _06754_ = sel_oi_one_hot_i[236] & i[192];
  assign _06755_ = sel_oi_one_hot_i[237] & i[208];
  assign _06756_ = _06755_ | _06754_;
  assign _06757_ = sel_oi_one_hot_i[238] & i[224];
  assign _06758_ = sel_oi_one_hot_i[239] & i[240];
  assign _06759_ = _06758_ | _06757_;
  assign _06760_ = _06759_ | _06756_;
  assign _06761_ = _06760_ | _06753_;
  assign o[224] = _06761_ | _06745_;
  assign _06763_ = i[7] & sel_oi_one_hot_i[16];
  assign _06764_ = i[23] & sel_oi_one_hot_i[17];
  assign _06765_ = _06764_ | _06763_;
  assign _06766_ = i[39] & sel_oi_one_hot_i[18];
  assign _06767_ = i[55] & sel_oi_one_hot_i[19];
  assign _06768_ = _06767_ | _06766_;
  assign _06769_ = _06768_ | _06765_;
  assign _06770_ = i[71] & sel_oi_one_hot_i[20];
  assign _06771_ = i[87] & sel_oi_one_hot_i[21];
  assign _06773_ = _06771_ | _06770_;
  assign _06774_ = i[103] & sel_oi_one_hot_i[22];
  assign _06775_ = i[119] & sel_oi_one_hot_i[23];
  assign _06776_ = _06775_ | _06774_;
  assign _06777_ = _06776_ | _06773_;
  assign _06778_ = _06777_ | _06769_;
  assign _06779_ = i[135] & sel_oi_one_hot_i[24];
  assign _06780_ = i[151] & sel_oi_one_hot_i[25];
  assign _06781_ = _06780_ | _06779_;
  assign _06782_ = i[167] & sel_oi_one_hot_i[26];
  assign _06784_ = i[183] & sel_oi_one_hot_i[27];
  assign _06785_ = _06784_ | _06782_;
  assign _06786_ = _06785_ | _06781_;
  assign _06787_ = i[199] & sel_oi_one_hot_i[28];
  assign _06788_ = i[215] & sel_oi_one_hot_i[29];
  assign _06789_ = _06788_ | _06787_;
  assign _06790_ = i[231] & sel_oi_one_hot_i[30];
  assign _06791_ = sel_oi_one_hot_i[31] & i[247];
  assign _06792_ = _06791_ | _06790_;
  assign _06793_ = _06792_ | _06789_;
  assign _06795_ = _06793_ | _06786_;
  assign o[23] = _06795_ | _06778_;
  assign _06796_ = sel_oi_one_hot_i[240] & i[15];
  assign _06797_ = sel_oi_one_hot_i[241] & i[31];
  assign _06798_ = _06797_ | _06796_;
  assign _06799_ = sel_oi_one_hot_i[242] & i[47];
  assign _06800_ = sel_oi_one_hot_i[243] & i[63];
  assign _06801_ = _06800_ | _06799_;
  assign _06802_ = _06801_ | _06798_;
  assign _06803_ = sel_oi_one_hot_i[244] & i[79];
  assign _06804_ = sel_oi_one_hot_i[245] & i[95];
  assign _06805_ = _06804_ | _06803_;
  assign _06806_ = sel_oi_one_hot_i[246] & i[111];
  assign _06807_ = sel_oi_one_hot_i[247] & i[127];
  assign _06808_ = _06807_ | _06806_;
  assign _06809_ = _06808_ | _06805_;
  assign _06810_ = _06809_ | _06802_;
  assign _06811_ = sel_oi_one_hot_i[248] & i[143];
  assign _06812_ = sel_oi_one_hot_i[249] & i[159];
  assign _06813_ = _06812_ | _06811_;
  assign _06815_ = sel_oi_one_hot_i[250] & i[175];
  assign _06816_ = sel_oi_one_hot_i[251] & i[191];
  assign _06817_ = _06816_ | _06815_;
  assign _06818_ = _06817_ | _06813_;
  assign _06819_ = sel_oi_one_hot_i[252] & i[207];
  assign _06820_ = sel_oi_one_hot_i[253] & i[223];
  assign _06821_ = _06820_ | _06819_;
  assign _06822_ = sel_oi_one_hot_i[254] & i[239];
  assign _06823_ = sel_oi_one_hot_i[255] & i[255];
  assign _06824_ = _06823_ | _06822_;
  assign _06826_ = _06824_ | _06821_;
  assign _06827_ = _06826_ | _06818_;
  assign o[255] = _06827_ | _06810_;
  assign _06828_ = sel_oi_one_hot_i[240] & i[14];
  assign _06829_ = sel_oi_one_hot_i[241] & i[30];
  assign _06830_ = _06829_ | _06828_;
  assign _06831_ = sel_oi_one_hot_i[242] & i[46];
  assign _06832_ = sel_oi_one_hot_i[243] & i[62];
  assign _06833_ = _06832_ | _06831_;
  assign _06834_ = _06833_ | _06830_;
  assign _06836_ = sel_oi_one_hot_i[244] & i[78];
  assign _06837_ = sel_oi_one_hot_i[245] & i[94];
  assign _06838_ = _06837_ | _06836_;
  assign _06839_ = sel_oi_one_hot_i[246] & i[110];
  assign _06840_ = sel_oi_one_hot_i[247] & i[126];
  assign _06841_ = _06840_ | _06839_;
  assign _06842_ = _06841_ | _06838_;
  assign _06843_ = _06842_ | _06834_;
  assign _06844_ = sel_oi_one_hot_i[248] & i[142];
  assign _06845_ = sel_oi_one_hot_i[249] & i[158];
  assign _06847_ = _06845_ | _06844_;
  assign _06848_ = sel_oi_one_hot_i[250] & i[174];
  assign _06849_ = sel_oi_one_hot_i[251] & i[190];
  assign _06850_ = _06849_ | _06848_;
  assign _06851_ = _06850_ | _06847_;
  assign _06852_ = sel_oi_one_hot_i[252] & i[206];
  assign _06853_ = sel_oi_one_hot_i[253] & i[222];
  assign _06854_ = _06853_ | _06852_;
  assign _06855_ = sel_oi_one_hot_i[254] & i[238];
  assign _06856_ = sel_oi_one_hot_i[255] & i[254];
  assign _06858_ = _06856_ | _06855_;
  assign _06859_ = _06858_ | _06854_;
  assign _06860_ = _06859_ | _06851_;
  assign o[254] = _06860_ | _06843_;
  assign _06861_ = sel_oi_one_hot_i[240] & i[13];
  assign _06862_ = sel_oi_one_hot_i[241] & i[29];
  assign _06863_ = _06862_ | _06861_;
  assign _06864_ = sel_oi_one_hot_i[242] & i[45];
  assign _06865_ = sel_oi_one_hot_i[243] & i[61];
  assign _06866_ = _06865_ | _06864_;
  assign _06868_ = _06866_ | _06863_;
  assign _06869_ = sel_oi_one_hot_i[244] & i[77];
  assign _06870_ = sel_oi_one_hot_i[245] & i[93];
  assign _06871_ = _06870_ | _06869_;
  assign _06872_ = sel_oi_one_hot_i[246] & i[109];
  assign _06873_ = sel_oi_one_hot_i[247] & i[125];
  assign _06874_ = _06873_ | _06872_;
  assign _06875_ = _06874_ | _06871_;
  assign _06876_ = _06875_ | _06868_;
  assign _06877_ = sel_oi_one_hot_i[248] & i[141];
  assign _06879_ = sel_oi_one_hot_i[249] & i[157];
  assign _06880_ = _06879_ | _06877_;
  assign _06881_ = sel_oi_one_hot_i[250] & i[173];
  assign _06882_ = sel_oi_one_hot_i[251] & i[189];
  assign _06883_ = _06882_ | _06881_;
  assign _06884_ = _06883_ | _06880_;
  assign _06885_ = sel_oi_one_hot_i[252] & i[205];
  assign _06886_ = sel_oi_one_hot_i[253] & i[221];
  assign _06887_ = _06886_ | _06885_;
  assign _06888_ = sel_oi_one_hot_i[254] & i[237];
  assign _06890_ = sel_oi_one_hot_i[255] & i[253];
  assign _06891_ = _06890_ | _06888_;
  assign _06892_ = _06891_ | _06887_;
  assign _06893_ = _06892_ | _06884_;
  assign o[253] = _06893_ | _06876_;
  assign _06894_ = sel_oi_one_hot_i[240] & i[12];
  assign _06895_ = sel_oi_one_hot_i[241] & i[28];
  assign _06896_ = _06895_ | _06894_;
  assign _06897_ = sel_oi_one_hot_i[242] & i[44];
  assign _06898_ = sel_oi_one_hot_i[243] & i[60];
  assign _06900_ = _06898_ | _06897_;
  assign _06901_ = _06900_ | _06896_;
  assign _06902_ = sel_oi_one_hot_i[244] & i[76];
  assign _06903_ = sel_oi_one_hot_i[245] & i[92];
  assign _06904_ = _06903_ | _06902_;
  assign _06905_ = sel_oi_one_hot_i[246] & i[108];
  assign _06906_ = sel_oi_one_hot_i[247] & i[124];
  assign _06907_ = _06906_ | _06905_;
  assign _06908_ = _06907_ | _06904_;
  assign _06909_ = _06908_ | _06901_;
  assign _06911_ = sel_oi_one_hot_i[248] & i[140];
  assign _06912_ = sel_oi_one_hot_i[249] & i[156];
  assign _06913_ = _06912_ | _06911_;
  assign _06914_ = sel_oi_one_hot_i[250] & i[172];
  assign _06915_ = sel_oi_one_hot_i[251] & i[188];
  assign _06916_ = _06915_ | _06914_;
  assign _06917_ = _06916_ | _06913_;
  assign _06918_ = sel_oi_one_hot_i[252] & i[204];
  assign _06919_ = sel_oi_one_hot_i[253] & i[220];
  assign _06920_ = _06919_ | _06918_;
  assign _06922_ = sel_oi_one_hot_i[254] & i[236];
  assign _06923_ = sel_oi_one_hot_i[255] & i[252];
  assign _06924_ = _06923_ | _06922_;
  assign _06925_ = _06924_ | _06920_;
  assign _06926_ = _06925_ | _06917_;
  assign o[252] = _06926_ | _06909_;
  assign _06927_ = i[6] & sel_oi_one_hot_i[16];
  assign _06928_ = i[22] & sel_oi_one_hot_i[17];
  assign _06929_ = _06928_ | _06927_;
  assign _06930_ = i[38] & sel_oi_one_hot_i[18];
  assign _06932_ = i[54] & sel_oi_one_hot_i[19];
  assign _06933_ = _06932_ | _06930_;
  assign _06934_ = _06933_ | _06929_;
  assign _06935_ = i[70] & sel_oi_one_hot_i[20];
  assign _06936_ = i[86] & sel_oi_one_hot_i[21];
  assign _06937_ = _06936_ | _06935_;
  assign _06938_ = i[102] & sel_oi_one_hot_i[22];
  assign _06939_ = i[118] & sel_oi_one_hot_i[23];
  assign _06940_ = _06939_ | _06938_;
  assign _06941_ = _06940_ | _06937_;
  assign _06943_ = _06941_ | _06934_;
  assign _06944_ = i[134] & sel_oi_one_hot_i[24];
  assign _06945_ = i[150] & sel_oi_one_hot_i[25];
  assign _06946_ = _06945_ | _06944_;
  assign _06947_ = i[166] & sel_oi_one_hot_i[26];
  assign _06948_ = i[182] & sel_oi_one_hot_i[27];
  assign _06949_ = _06948_ | _06947_;
  assign _06950_ = _06949_ | _06946_;
  assign _06951_ = i[198] & sel_oi_one_hot_i[28];
  assign _06952_ = i[214] & sel_oi_one_hot_i[29];
  assign _06954_ = _06952_ | _06951_;
  assign _06955_ = i[230] & sel_oi_one_hot_i[30];
  assign _06956_ = sel_oi_one_hot_i[31] & i[246];
  assign _06957_ = _06956_ | _06955_;
  assign _06958_ = _06957_ | _06954_;
  assign _06959_ = _06958_ | _06950_;
  assign o[22] = _06959_ | _06943_;
  assign _06960_ = sel_oi_one_hot_i[240] & i[11];
  assign _06961_ = sel_oi_one_hot_i[241] & i[27];
  assign _06962_ = _06961_ | _06960_;
  assign _06964_ = sel_oi_one_hot_i[242] & i[43];
  assign _06965_ = sel_oi_one_hot_i[243] & i[59];
  assign _06966_ = _06965_ | _06964_;
  assign _06967_ = _06966_ | _06962_;
  assign _06968_ = sel_oi_one_hot_i[244] & i[75];
  assign _06969_ = sel_oi_one_hot_i[245] & i[91];
  assign _06970_ = _06969_ | _06968_;
  assign _06971_ = sel_oi_one_hot_i[246] & i[107];
  assign _06972_ = sel_oi_one_hot_i[247] & i[123];
  assign _06973_ = _06972_ | _06971_;
  assign _06975_ = _06973_ | _06970_;
  assign _06976_ = _06975_ | _06967_;
  assign _06977_ = sel_oi_one_hot_i[248] & i[139];
  assign _06978_ = sel_oi_one_hot_i[249] & i[155];
  assign _06979_ = _06978_ | _06977_;
  assign _06980_ = sel_oi_one_hot_i[250] & i[171];
  assign _06981_ = sel_oi_one_hot_i[251] & i[187];
  assign _06982_ = _06981_ | _06980_;
  assign _06983_ = _06982_ | _06979_;
  assign _06984_ = sel_oi_one_hot_i[252] & i[203];
  assign _06986_ = sel_oi_one_hot_i[253] & i[219];
  assign _06987_ = _06986_ | _06984_;
  assign _06988_ = sel_oi_one_hot_i[254] & i[235];
  assign _06989_ = sel_oi_one_hot_i[255] & i[251];
  assign _06990_ = _06989_ | _06988_;
  assign _06991_ = _06990_ | _06987_;
  assign _06992_ = _06991_ | _06983_;
  assign o[251] = _06992_ | _06976_;
  assign _06993_ = sel_oi_one_hot_i[240] & i[10];
  assign _06994_ = sel_oi_one_hot_i[241] & i[26];
  assign _06996_ = _06994_ | _06993_;
  assign _06997_ = sel_oi_one_hot_i[242] & i[42];
  assign _06998_ = sel_oi_one_hot_i[243] & i[58];
  assign _06999_ = _06998_ | _06997_;
  assign _07000_ = _06999_ | _06996_;
  assign _07001_ = sel_oi_one_hot_i[244] & i[74];
  assign _07002_ = sel_oi_one_hot_i[245] & i[90];
  assign _07003_ = _07002_ | _07001_;
  assign _07004_ = sel_oi_one_hot_i[246] & i[106];
  assign _07005_ = sel_oi_one_hot_i[247] & i[122];
  assign _07007_ = _07005_ | _07004_;
  assign _07008_ = _07007_ | _07003_;
  assign _07009_ = _07008_ | _07000_;
  assign _07010_ = sel_oi_one_hot_i[248] & i[138];
  assign _07011_ = sel_oi_one_hot_i[249] & i[154];
  assign _07012_ = _07011_ | _07010_;
  assign _07013_ = sel_oi_one_hot_i[250] & i[170];
  assign _07014_ = sel_oi_one_hot_i[251] & i[186];
  assign _07015_ = _07014_ | _07013_;
  assign _07016_ = _07015_ | _07012_;
  assign _07018_ = sel_oi_one_hot_i[252] & i[202];
  assign _07019_ = sel_oi_one_hot_i[253] & i[218];
  assign _07020_ = _07019_ | _07018_;
  assign _07021_ = sel_oi_one_hot_i[254] & i[234];
  assign _07022_ = sel_oi_one_hot_i[255] & i[250];
  assign _07023_ = _07022_ | _07021_;
  assign _07024_ = _07023_ | _07020_;
  assign _07025_ = _07024_ | _07016_;
  assign o[250] = _07025_ | _07009_;
  assign _07026_ = sel_oi_one_hot_i[240] & i[9];
  assign _07028_ = sel_oi_one_hot_i[241] & i[25];
  assign _07029_ = _07028_ | _07026_;
  assign _07030_ = sel_oi_one_hot_i[242] & i[41];
  assign _07031_ = sel_oi_one_hot_i[243] & i[57];
  assign _07032_ = _07031_ | _07030_;
  assign _07033_ = _07032_ | _07029_;
  assign _07034_ = sel_oi_one_hot_i[244] & i[73];
  assign _07035_ = sel_oi_one_hot_i[245] & i[89];
  assign _07036_ = _07035_ | _07034_;
  assign _07037_ = sel_oi_one_hot_i[246] & i[105];
  assign _07039_ = sel_oi_one_hot_i[247] & i[121];
  assign _07040_ = _07039_ | _07037_;
  assign _07041_ = _07040_ | _07036_;
  assign _07042_ = _07041_ | _07033_;
  assign _07043_ = sel_oi_one_hot_i[248] & i[137];
  assign _07044_ = sel_oi_one_hot_i[249] & i[153];
  assign _07045_ = _07044_ | _07043_;
  assign _07046_ = sel_oi_one_hot_i[250] & i[169];
  assign _07047_ = sel_oi_one_hot_i[251] & i[185];
  assign _07048_ = _07047_ | _07046_;
  assign _07050_ = _07048_ | _07045_;
  assign _07051_ = sel_oi_one_hot_i[252] & i[201];
  assign _07052_ = sel_oi_one_hot_i[253] & i[217];
  assign _07053_ = _07052_ | _07051_;
  assign _07054_ = sel_oi_one_hot_i[254] & i[233];
  assign _07055_ = sel_oi_one_hot_i[255] & i[249];
  assign _07056_ = _07055_ | _07054_;
  assign _07057_ = _07056_ | _07053_;
  assign _07058_ = _07057_ | _07050_;
  assign o[249] = _07058_ | _07042_;
  assign _07060_ = sel_oi_one_hot_i[240] & i[8];
  assign _07061_ = sel_oi_one_hot_i[241] & i[24];
  assign _07062_ = _07061_ | _07060_;
  assign _07063_ = sel_oi_one_hot_i[242] & i[40];
  assign _07064_ = sel_oi_one_hot_i[243] & i[56];
  assign _07065_ = _07064_ | _07063_;
  assign _07066_ = _07065_ | _07062_;
  assign _07067_ = sel_oi_one_hot_i[244] & i[72];
  assign _07068_ = sel_oi_one_hot_i[245] & i[88];
  assign _07069_ = _07068_ | _07067_;
  assign _07071_ = sel_oi_one_hot_i[246] & i[104];
  assign _07072_ = sel_oi_one_hot_i[247] & i[120];
  assign _07073_ = _07072_ | _07071_;
  assign _07074_ = _07073_ | _07069_;
  assign _07075_ = _07074_ | _07066_;
  assign _07076_ = sel_oi_one_hot_i[248] & i[136];
  assign _07077_ = sel_oi_one_hot_i[249] & i[152];
  assign _07078_ = _07077_ | _07076_;
  assign _07079_ = sel_oi_one_hot_i[250] & i[168];
  assign _07080_ = sel_oi_one_hot_i[251] & i[184];
  assign _07082_ = _07080_ | _07079_;
  assign _07083_ = _07082_ | _07078_;
  assign _07084_ = sel_oi_one_hot_i[252] & i[200];
  assign _07085_ = sel_oi_one_hot_i[253] & i[216];
  assign _07086_ = _07085_ | _07084_;
  assign _07087_ = sel_oi_one_hot_i[254] & i[232];
  assign _07088_ = sel_oi_one_hot_i[255] & i[248];
  assign _07089_ = _07088_ | _07087_;
  assign _07090_ = _07089_ | _07086_;
  assign _07091_ = _07090_ | _07083_;
  assign o[248] = _07091_ | _07075_;
  assign _07093_ = sel_oi_one_hot_i[240] & i[7];
  assign _07094_ = sel_oi_one_hot_i[241] & i[23];
  assign _07095_ = _07094_ | _07093_;
  assign _07096_ = sel_oi_one_hot_i[242] & i[39];
  assign _07097_ = sel_oi_one_hot_i[243] & i[55];
  assign _07098_ = _07097_ | _07096_;
  assign _07099_ = _07098_ | _07095_;
  assign _07100_ = sel_oi_one_hot_i[244] & i[71];
  assign _07101_ = sel_oi_one_hot_i[245] & i[87];
  assign _07103_ = _07101_ | _07100_;
  assign _07104_ = sel_oi_one_hot_i[246] & i[103];
  assign _07105_ = sel_oi_one_hot_i[247] & i[119];
  assign _07106_ = _07105_ | _07104_;
  assign _07107_ = _07106_ | _07103_;
  assign _07108_ = _07107_ | _07099_;
  assign _07109_ = sel_oi_one_hot_i[248] & i[135];
  assign _07110_ = sel_oi_one_hot_i[249] & i[151];
  assign _07111_ = _07110_ | _07109_;
  assign _07112_ = sel_oi_one_hot_i[250] & i[167];
  assign _07114_ = sel_oi_one_hot_i[251] & i[183];
  assign _07115_ = _07114_ | _07112_;
  assign _07116_ = _07115_ | _07111_;
  assign _07117_ = sel_oi_one_hot_i[252] & i[199];
  assign _07118_ = sel_oi_one_hot_i[253] & i[215];
  assign _07119_ = _07118_ | _07117_;
  assign _07120_ = sel_oi_one_hot_i[254] & i[231];
  assign _07121_ = sel_oi_one_hot_i[255] & i[247];
  assign _07122_ = _07121_ | _07120_;
  assign _07123_ = _07122_ | _07119_;
  assign _07125_ = _07123_ | _07116_;
  assign o[247] = _07125_ | _07108_;
  assign _07126_ = sel_oi_one_hot_i[240] & i[6];
  assign _07127_ = sel_oi_one_hot_i[241] & i[22];
  assign _07128_ = _07127_ | _07126_;
  assign _07129_ = sel_oi_one_hot_i[242] & i[38];
  assign _07130_ = sel_oi_one_hot_i[243] & i[54];
  assign _07131_ = _07130_ | _07129_;
  assign _07132_ = _07131_ | _07128_;
  assign _07133_ = sel_oi_one_hot_i[244] & i[70];
  assign _07134_ = sel_oi_one_hot_i[245] & i[86];
  assign _07135_ = _07134_ | _07133_;
  assign _07136_ = sel_oi_one_hot_i[246] & i[102];
  assign _07137_ = sel_oi_one_hot_i[247] & i[118];
  assign _07138_ = _07137_ | _07136_;
  assign _07139_ = _07138_ | _07135_;
  assign _07140_ = _07139_ | _07132_;
  assign _07141_ = sel_oi_one_hot_i[248] & i[134];
  assign _07142_ = sel_oi_one_hot_i[249] & i[150];
  assign _07143_ = _07142_ | _07141_;
  assign _07145_ = sel_oi_one_hot_i[250] & i[166];
  assign _07146_ = sel_oi_one_hot_i[251] & i[182];
  assign _07147_ = _07146_ | _07145_;
  assign _07148_ = _07147_ | _07143_;
  assign _07149_ = sel_oi_one_hot_i[252] & i[198];
  assign _07150_ = sel_oi_one_hot_i[253] & i[214];
  assign _07151_ = _07150_ | _07149_;
  assign _07152_ = sel_oi_one_hot_i[254] & i[230];
  assign _07153_ = sel_oi_one_hot_i[255] & i[246];
  assign _07154_ = _07153_ | _07152_;
  assign _07156_ = _07154_ | _07151_;
  assign _07157_ = _07156_ | _07148_;
  assign o[246] = _07157_ | _07140_;
  assign _07158_ = sel_oi_one_hot_i[240] & i[5];
  assign _07159_ = sel_oi_one_hot_i[241] & i[21];
  assign _07160_ = _07159_ | _07158_;
  assign _07161_ = sel_oi_one_hot_i[242] & i[37];
  assign _07162_ = sel_oi_one_hot_i[243] & i[53];
  assign _07163_ = _07162_ | _07161_;
  assign _07164_ = _07163_ | _07160_;
  assign _07166_ = sel_oi_one_hot_i[244] & i[69];
  assign _07167_ = sel_oi_one_hot_i[245] & i[85];
  assign _07168_ = _07167_ | _07166_;
  assign _07169_ = sel_oi_one_hot_i[246] & i[101];
  assign _07170_ = sel_oi_one_hot_i[247] & i[117];
  assign _07171_ = _07170_ | _07169_;
  assign _07172_ = _07171_ | _07168_;
  assign _07173_ = _07172_ | _07164_;
  assign _07174_ = sel_oi_one_hot_i[248] & i[133];
  assign _07175_ = sel_oi_one_hot_i[249] & i[149];
  assign _07177_ = _07175_ | _07174_;
  assign _07178_ = sel_oi_one_hot_i[250] & i[165];
  assign _07179_ = sel_oi_one_hot_i[251] & i[181];
  assign _07180_ = _07179_ | _07178_;
  assign _07181_ = _07180_ | _07177_;
  assign _07182_ = sel_oi_one_hot_i[252] & i[197];
  assign _07183_ = sel_oi_one_hot_i[253] & i[213];
  assign _07184_ = _07183_ | _07182_;
  assign _07185_ = sel_oi_one_hot_i[254] & i[229];
  assign _07186_ = sel_oi_one_hot_i[255] & i[245];
  assign _07188_ = _07186_ | _07185_;
  assign _07189_ = _07188_ | _07184_;
  assign _07190_ = _07189_ | _07181_;
  assign o[245] = _07190_ | _07173_;
  assign _07191_ = sel_oi_one_hot_i[240] & i[4];
  assign _07192_ = sel_oi_one_hot_i[241] & i[20];
  assign _07193_ = _07192_ | _07191_;
  assign _07194_ = sel_oi_one_hot_i[242] & i[36];
  assign _07195_ = sel_oi_one_hot_i[243] & i[52];
  assign _07196_ = _07195_ | _07194_;
  assign _07198_ = _07196_ | _07193_;
  assign _07199_ = sel_oi_one_hot_i[244] & i[68];
  assign _07200_ = sel_oi_one_hot_i[245] & i[84];
  assign _07201_ = _07200_ | _07199_;
  assign _07202_ = sel_oi_one_hot_i[246] & i[100];
  assign _07203_ = sel_oi_one_hot_i[247] & i[116];
  assign _07204_ = _07203_ | _07202_;
  assign _07205_ = _07204_ | _07201_;
  assign _07206_ = _07205_ | _07198_;
  assign _07207_ = sel_oi_one_hot_i[248] & i[132];
  assign _07209_ = sel_oi_one_hot_i[249] & i[148];
  assign _07210_ = _07209_ | _07207_;
  assign _07211_ = sel_oi_one_hot_i[250] & i[164];
  assign _07212_ = sel_oi_one_hot_i[251] & i[180];
  assign _07213_ = _07212_ | _07211_;
  assign _07214_ = _07213_ | _07210_;
  assign _07215_ = sel_oi_one_hot_i[252] & i[196];
  assign _07216_ = sel_oi_one_hot_i[253] & i[212];
  assign _07217_ = _07216_ | _07215_;
  assign _07218_ = sel_oi_one_hot_i[254] & i[228];
  assign _07220_ = sel_oi_one_hot_i[255] & i[244];
  assign _07221_ = _07220_ | _07218_;
  assign _07222_ = _07221_ | _07217_;
  assign _07223_ = _07222_ | _07214_;
  assign o[244] = _07223_ | _07206_;
  assign _07224_ = sel_oi_one_hot_i[240] & i[3];
  assign _07225_ = sel_oi_one_hot_i[241] & i[19];
  assign _07226_ = _07225_ | _07224_;
  assign _07227_ = sel_oi_one_hot_i[242] & i[35];
  assign _07228_ = sel_oi_one_hot_i[243] & i[51];
  assign _07230_ = _07228_ | _07227_;
  assign _07231_ = _07230_ | _07226_;
  assign _07232_ = sel_oi_one_hot_i[244] & i[67];
  assign _07233_ = sel_oi_one_hot_i[245] & i[83];
  assign _07234_ = _07233_ | _07232_;
  assign _07235_ = sel_oi_one_hot_i[246] & i[99];
  assign _07236_ = sel_oi_one_hot_i[247] & i[115];
  assign _07237_ = _07236_ | _07235_;
  assign _07238_ = _07237_ | _07234_;
  assign _07239_ = _07238_ | _07231_;
  assign _07241_ = sel_oi_one_hot_i[248] & i[131];
  assign _07242_ = sel_oi_one_hot_i[249] & i[147];
  assign _07243_ = _07242_ | _07241_;
  assign _07244_ = sel_oi_one_hot_i[250] & i[163];
  assign _07245_ = sel_oi_one_hot_i[251] & i[179];
  assign _07246_ = _07245_ | _07244_;
  assign _07247_ = _07246_ | _07243_;
  assign _07248_ = sel_oi_one_hot_i[252] & i[195];
  assign _07249_ = sel_oi_one_hot_i[253] & i[211];
  assign _07250_ = _07249_ | _07248_;
  assign _07252_ = sel_oi_one_hot_i[254] & i[227];
  assign _07253_ = sel_oi_one_hot_i[255] & i[243];
  assign _07254_ = _07253_ | _07252_;
  assign _07255_ = _07254_ | _07250_;
  assign _07256_ = _07255_ | _07247_;
  assign o[243] = _07256_ | _07239_;
  assign _07257_ = sel_oi_one_hot_i[240] & i[2];
  assign _07258_ = sel_oi_one_hot_i[241] & i[18];
  assign _07259_ = _07258_ | _07257_;
  assign _07260_ = sel_oi_one_hot_i[242] & i[34];
  assign _07262_ = sel_oi_one_hot_i[243] & i[50];
  assign _07263_ = _07262_ | _07260_;
  assign _07264_ = _07263_ | _07259_;
  assign _07265_ = sel_oi_one_hot_i[244] & i[66];
  assign _07266_ = sel_oi_one_hot_i[245] & i[82];
  assign _07267_ = _07266_ | _07265_;
  assign _07268_ = sel_oi_one_hot_i[246] & i[98];
  assign _07269_ = sel_oi_one_hot_i[247] & i[114];
  assign _07270_ = _07269_ | _07268_;
  assign _07271_ = _07270_ | _07267_;
  assign _07273_ = _07271_ | _07264_;
  assign _07274_ = sel_oi_one_hot_i[248] & i[130];
  assign _07275_ = sel_oi_one_hot_i[249] & i[146];
  assign _07276_ = _07275_ | _07274_;
  assign _07277_ = sel_oi_one_hot_i[250] & i[162];
  assign _07278_ = sel_oi_one_hot_i[251] & i[178];
  assign _07279_ = _07278_ | _07277_;
  assign _07280_ = _07279_ | _07276_;
  assign _07281_ = sel_oi_one_hot_i[252] & i[194];
  assign _07282_ = sel_oi_one_hot_i[253] & i[210];
  assign _07284_ = _07282_ | _07281_;
  assign _07285_ = sel_oi_one_hot_i[254] & i[226];
  assign _07286_ = sel_oi_one_hot_i[255] & i[242];
  assign _07287_ = _07286_ | _07285_;
  assign _07288_ = _07287_ | _07284_;
  assign _07289_ = _07288_ | _07280_;
  assign o[242] = _07289_ | _07273_;
  assign _07290_ = i[5] & sel_oi_one_hot_i[16];
  assign _07291_ = i[21] & sel_oi_one_hot_i[17];
  assign _07292_ = _07291_ | _07290_;
  assign _07294_ = i[37] & sel_oi_one_hot_i[18];
  assign _07295_ = i[53] & sel_oi_one_hot_i[19];
  assign _07296_ = _07295_ | _07294_;
  assign _07297_ = _07296_ | _07292_;
  assign _07298_ = i[69] & sel_oi_one_hot_i[20];
  assign _07299_ = i[85] & sel_oi_one_hot_i[21];
  assign _07300_ = _07299_ | _07298_;
  assign _07301_ = i[101] & sel_oi_one_hot_i[22];
  assign _07302_ = i[117] & sel_oi_one_hot_i[23];
  assign _07303_ = _07302_ | _07301_;
  assign _07305_ = _07303_ | _07300_;
  assign _07306_ = _07305_ | _07297_;
  assign _07307_ = i[133] & sel_oi_one_hot_i[24];
  assign _07308_ = i[149] & sel_oi_one_hot_i[25];
  assign _07309_ = _07308_ | _07307_;
  assign _07310_ = i[165] & sel_oi_one_hot_i[26];
  assign _07311_ = i[181] & sel_oi_one_hot_i[27];
  assign _07312_ = _07311_ | _07310_;
  assign _07313_ = _07312_ | _07309_;
  assign _07314_ = i[197] & sel_oi_one_hot_i[28];
  assign _07316_ = i[213] & sel_oi_one_hot_i[29];
  assign _07317_ = _07316_ | _07314_;
  assign _07318_ = i[229] & sel_oi_one_hot_i[30];
  assign _07319_ = sel_oi_one_hot_i[31] & i[245];
  assign _07320_ = _07319_ | _07318_;
  assign _07321_ = _07320_ | _07317_;
  assign _07322_ = _07321_ | _07313_;
  assign o[21] = _07322_ | _07306_;
  assign _07323_ = sel_oi_one_hot_i[240] & i[1];
  assign _07324_ = sel_oi_one_hot_i[241] & i[17];
  assign _07326_ = _07324_ | _07323_;
  assign _07327_ = sel_oi_one_hot_i[242] & i[33];
  assign _07328_ = sel_oi_one_hot_i[243] & i[49];
  assign _07329_ = _07328_ | _07327_;
  assign _07330_ = _07329_ | _07326_;
  assign _07331_ = sel_oi_one_hot_i[244] & i[65];
  assign _07332_ = sel_oi_one_hot_i[245] & i[81];
  assign _07333_ = _07332_ | _07331_;
  assign _07334_ = sel_oi_one_hot_i[246] & i[97];
  assign _07335_ = sel_oi_one_hot_i[247] & i[113];
  assign _07337_ = _07335_ | _07334_;
  assign _07338_ = _07337_ | _07333_;
  assign _07339_ = _07338_ | _07330_;
  assign _07340_ = sel_oi_one_hot_i[248] & i[129];
  assign _07341_ = sel_oi_one_hot_i[249] & i[145];
  assign _07342_ = _07341_ | _07340_;
  assign _07343_ = sel_oi_one_hot_i[250] & i[161];
  assign _07344_ = sel_oi_one_hot_i[251] & i[177];
  assign _07345_ = _07344_ | _07343_;
  assign _07346_ = _07345_ | _07342_;
  assign _07348_ = sel_oi_one_hot_i[252] & i[193];
  assign _07349_ = sel_oi_one_hot_i[253] & i[209];
  assign _07350_ = _07349_ | _07348_;
  assign _07351_ = sel_oi_one_hot_i[254] & i[225];
  assign _07352_ = sel_oi_one_hot_i[255] & i[241];
  assign _07353_ = _07352_ | _07351_;
  assign _07354_ = _07353_ | _07350_;
  assign _07355_ = _07354_ | _07346_;
  assign o[241] = _07355_ | _07339_;
  assign _07356_ = sel_oi_one_hot_i[240] & i[0];
  assign _07358_ = sel_oi_one_hot_i[241] & i[16];
  assign _07359_ = _07358_ | _07356_;
  assign _07360_ = sel_oi_one_hot_i[242] & i[32];
  assign _07361_ = sel_oi_one_hot_i[243] & i[48];
  assign _07362_ = _07361_ | _07360_;
  assign _07363_ = _07362_ | _07359_;
  assign _07364_ = sel_oi_one_hot_i[244] & i[64];
  assign _07365_ = sel_oi_one_hot_i[245] & i[80];
  assign _07366_ = _07365_ | _07364_;
  assign _07367_ = sel_oi_one_hot_i[246] & i[96];
  assign _07369_ = sel_oi_one_hot_i[247] & i[112];
  assign _07370_ = _07369_ | _07367_;
  assign _07371_ = _07370_ | _07366_;
  assign _07372_ = _07371_ | _07363_;
  assign _07373_ = sel_oi_one_hot_i[248] & i[128];
  assign _07374_ = sel_oi_one_hot_i[249] & i[144];
  assign _07375_ = _07374_ | _07373_;
  assign _07376_ = sel_oi_one_hot_i[250] & i[160];
  assign _07377_ = sel_oi_one_hot_i[251] & i[176];
  assign _07378_ = _07377_ | _07376_;
  assign _07380_ = _07378_ | _07375_;
  assign _07381_ = sel_oi_one_hot_i[252] & i[192];
  assign _07382_ = sel_oi_one_hot_i[253] & i[208];
  assign _07383_ = _07382_ | _07381_;
  assign _07384_ = sel_oi_one_hot_i[254] & i[224];
  assign _07385_ = sel_oi_one_hot_i[255] & i[240];
  assign _07386_ = _07385_ | _07384_;
  assign _07387_ = _07386_ | _07383_;
  assign _07388_ = _07387_ | _07380_;
  assign o[240] = _07388_ | _07372_;
  assign _07390_ = i[4] & sel_oi_one_hot_i[16];
  assign _07391_ = i[20] & sel_oi_one_hot_i[17];
  assign _07392_ = _07391_ | _07390_;
  assign _07393_ = i[36] & sel_oi_one_hot_i[18];
  assign _07394_ = i[52] & sel_oi_one_hot_i[19];
  assign _07395_ = _07394_ | _07393_;
  assign _07396_ = _07395_ | _07392_;
  assign _07397_ = i[68] & sel_oi_one_hot_i[20];
  assign _07398_ = i[84] & sel_oi_one_hot_i[21];
  assign _07399_ = _07398_ | _07397_;
  assign _07401_ = i[100] & sel_oi_one_hot_i[22];
  assign _07402_ = i[116] & sel_oi_one_hot_i[23];
  assign _07403_ = _07402_ | _07401_;
  assign _07404_ = _07403_ | _07399_;
  assign _07405_ = _07404_ | _07396_;
  assign _07406_ = i[132] & sel_oi_one_hot_i[24];
  assign _07407_ = i[148] & sel_oi_one_hot_i[25];
  assign _07408_ = _07407_ | _07406_;
  assign _07409_ = i[164] & sel_oi_one_hot_i[26];
  assign _07410_ = i[180] & sel_oi_one_hot_i[27];
  assign _07412_ = _07410_ | _07409_;
  assign _07413_ = _07412_ | _07408_;
  assign _07414_ = i[196] & sel_oi_one_hot_i[28];
  assign _07415_ = i[212] & sel_oi_one_hot_i[29];
  assign _07416_ = _07415_ | _07414_;
  assign _07417_ = i[228] & sel_oi_one_hot_i[30];
  assign _07418_ = sel_oi_one_hot_i[31] & i[244];
  assign _07419_ = _07418_ | _07417_;
  assign _07420_ = _07419_ | _07416_;
  assign _07421_ = _07420_ | _07413_;
  assign o[20] = _07421_ | _07405_;
  assign _07423_ = i[3] & sel_oi_one_hot_i[16];
  assign _07424_ = i[19] & sel_oi_one_hot_i[17];
  assign _07425_ = _07424_ | _07423_;
  assign _07426_ = i[35] & sel_oi_one_hot_i[18];
  assign _07427_ = i[51] & sel_oi_one_hot_i[19];
  assign _07428_ = _07427_ | _07426_;
  assign _07429_ = _07428_ | _07425_;
  assign _07430_ = i[67] & sel_oi_one_hot_i[20];
  assign _07431_ = i[83] & sel_oi_one_hot_i[21];
  assign _07433_ = _07431_ | _07430_;
  assign _07434_ = i[99] & sel_oi_one_hot_i[22];
  assign _07435_ = i[115] & sel_oi_one_hot_i[23];
  assign _07436_ = _07435_ | _07434_;
  assign _07437_ = _07436_ | _07433_;
  assign _07438_ = _07437_ | _07429_;
  assign _07439_ = i[131] & sel_oi_one_hot_i[24];
  assign _07440_ = i[147] & sel_oi_one_hot_i[25];
  assign _07441_ = _07440_ | _07439_;
  assign _07442_ = i[163] & sel_oi_one_hot_i[26];
  assign _07444_ = i[179] & sel_oi_one_hot_i[27];
  assign _07445_ = _07444_ | _07442_;
  assign _07446_ = _07445_ | _07441_;
  assign _07447_ = i[195] & sel_oi_one_hot_i[28];
  assign _07448_ = i[211] & sel_oi_one_hot_i[29];
  assign _07449_ = _07448_ | _07447_;
  assign _07450_ = i[227] & sel_oi_one_hot_i[30];
  assign _07451_ = sel_oi_one_hot_i[31] & i[243];
  assign _07452_ = _07451_ | _07450_;
  assign _07453_ = _07452_ | _07449_;
  assign _07455_ = _07453_ | _07446_;
  assign o[19] = _07455_ | _07438_;
  assign _07456_ = i[2] & sel_oi_one_hot_i[16];
  assign _07457_ = i[18] & sel_oi_one_hot_i[17];
  assign _07458_ = _07457_ | _07456_;
  assign _07459_ = i[34] & sel_oi_one_hot_i[18];
  assign _07460_ = i[50] & sel_oi_one_hot_i[19];
  assign _07461_ = _07460_ | _07459_;
  assign _07462_ = _07461_ | _07458_;
  assign _07463_ = i[66] & sel_oi_one_hot_i[20];
  assign _07464_ = i[82] & sel_oi_one_hot_i[21];
  assign _07465_ = _07464_ | _07463_;
  assign _07466_ = i[98] & sel_oi_one_hot_i[22];
  assign _07467_ = i[114] & sel_oi_one_hot_i[23];
  assign _07468_ = _07467_ | _07466_;
  assign _07469_ = _07468_ | _07465_;
  assign _07470_ = _07469_ | _07462_;
  assign _07471_ = i[130] & sel_oi_one_hot_i[24];
  assign _07472_ = i[146] & sel_oi_one_hot_i[25];
  assign _07473_ = _07472_ | _07471_;
  assign _07475_ = i[162] & sel_oi_one_hot_i[26];
  assign _07476_ = i[178] & sel_oi_one_hot_i[27];
  assign _07477_ = _07476_ | _07475_;
  assign _07478_ = _07477_ | _07473_;
  assign _07479_ = i[194] & sel_oi_one_hot_i[28];
  assign _07480_ = i[210] & sel_oi_one_hot_i[29];
  assign _07481_ = _07480_ | _07479_;
  assign _07482_ = i[226] & sel_oi_one_hot_i[30];
  assign _07483_ = sel_oi_one_hot_i[31] & i[242];
  assign _07484_ = _07483_ | _07482_;
  assign _07486_ = _07484_ | _07481_;
  assign _07487_ = _07486_ | _07478_;
  assign o[18] = _07487_ | _07470_;
  assign _07488_ = i[1] & sel_oi_one_hot_i[16];
  assign _07489_ = i[17] & sel_oi_one_hot_i[17];
  assign _07490_ = _07489_ | _07488_;
  assign _07491_ = i[33] & sel_oi_one_hot_i[18];
  assign _07492_ = i[49] & sel_oi_one_hot_i[19];
  assign _07493_ = _07492_ | _07491_;
  assign _07494_ = _07493_ | _07490_;
  assign _07496_ = i[65] & sel_oi_one_hot_i[20];
  assign _07497_ = i[81] & sel_oi_one_hot_i[21];
  assign _07498_ = _07497_ | _07496_;
  assign _07499_ = i[97] & sel_oi_one_hot_i[22];
  assign _07500_ = i[113] & sel_oi_one_hot_i[23];
  assign _07501_ = _07500_ | _07499_;
  assign _07502_ = _07501_ | _07498_;
  assign _07503_ = _07502_ | _07494_;
  assign _07504_ = i[129] & sel_oi_one_hot_i[24];
  assign _07505_ = i[145] & sel_oi_one_hot_i[25];
  assign _07507_ = _07505_ | _07504_;
  assign _07508_ = i[161] & sel_oi_one_hot_i[26];
  assign _07509_ = i[177] & sel_oi_one_hot_i[27];
  assign _07510_ = _07509_ | _07508_;
  assign _07511_ = _07510_ | _07507_;
  assign _07512_ = i[193] & sel_oi_one_hot_i[28];
  assign _07513_ = i[209] & sel_oi_one_hot_i[29];
  assign _07514_ = _07513_ | _07512_;
  assign _07515_ = i[225] & sel_oi_one_hot_i[30];
  assign _07516_ = sel_oi_one_hot_i[31] & i[241];
  assign _07518_ = _07516_ | _07515_;
  assign _07519_ = _07518_ | _07514_;
  assign _07520_ = _07519_ | _07511_;
  assign o[17] = _07520_ | _07503_;
  assign _07521_ = sel_oi_one_hot_i[16] & i[0];
  assign _07522_ = sel_oi_one_hot_i[17] & i[16];
  assign _07523_ = _07522_ | _07521_;
  assign _07524_ = sel_oi_one_hot_i[18] & i[32];
  assign _07525_ = sel_oi_one_hot_i[19] & i[48];
  assign _07526_ = _07525_ | _07524_;
  assign _07528_ = _07526_ | _07523_;
  assign _07529_ = sel_oi_one_hot_i[20] & i[64];
  assign _07530_ = sel_oi_one_hot_i[21] & i[80];
  assign _07531_ = _07530_ | _07529_;
  assign _07532_ = sel_oi_one_hot_i[22] & i[96];
  assign _07533_ = sel_oi_one_hot_i[23] & i[112];
  assign _07534_ = _07533_ | _07532_;
  assign _07535_ = _07534_ | _07531_;
  assign _07536_ = _07535_ | _07528_;
  assign _07537_ = sel_oi_one_hot_i[24] & i[128];
  assign _07539_ = sel_oi_one_hot_i[25] & i[144];
  assign _07540_ = _07539_ | _07537_;
  assign _07541_ = sel_oi_one_hot_i[26] & i[160];
  assign _07542_ = sel_oi_one_hot_i[27] & i[176];
  assign _07543_ = _07542_ | _07541_;
  assign _07544_ = _07543_ | _07540_;
  assign _07545_ = sel_oi_one_hot_i[28] & i[192];
  assign _07546_ = sel_oi_one_hot_i[29] & i[208];
  assign _07547_ = _07546_ | _07545_;
  assign _07548_ = i[224] & sel_oi_one_hot_i[30];
  assign _07550_ = sel_oi_one_hot_i[31] & i[240];
  assign _07551_ = _07550_ | _07548_;
  assign _07552_ = _07551_ | _07547_;
  assign _07553_ = _07552_ | _07544_;
  assign o[16] = _07553_ | _07536_;
  assign _06484_ = sel_oi_one_hot_i[32] & i[15];
  assign _06495_ = sel_oi_one_hot_i[33] & i[31];
  assign _06505_ = _06495_ | _06484_;
  assign _06516_ = sel_oi_one_hot_i[34] & i[47];
  assign _06527_ = sel_oi_one_hot_i[35] & i[63];
  assign _06537_ = _06527_ | _06516_;
  assign _06548_ = _06537_ | _06505_;
  assign _06559_ = sel_oi_one_hot_i[36] & i[79];
  assign _06569_ = sel_oi_one_hot_i[37] & i[95];
  assign _06580_ = _06569_ | _06559_;
  assign _06591_ = sel_oi_one_hot_i[38] & i[111];
  assign _06601_ = sel_oi_one_hot_i[39] & i[127];
  assign _06612_ = _06601_ | _06591_;
  assign _06623_ = _06612_ | _06580_;
  assign _06633_ = _06623_ | _06548_;
  assign _06644_ = sel_oi_one_hot_i[40] & i[143];
  assign _06655_ = sel_oi_one_hot_i[41] & i[159];
  assign _06665_ = _06655_ | _06644_;
  assign _06676_ = sel_oi_one_hot_i[42] & i[175];
  assign _06687_ = sel_oi_one_hot_i[43] & i[191];
  assign _06697_ = _06687_ | _06676_;
  assign _06708_ = _06697_ | _06665_;
  assign _06719_ = sel_oi_one_hot_i[44] & i[207];
  assign _06729_ = sel_oi_one_hot_i[45] & i[223];
  assign _06740_ = _06729_ | _06719_;
  assign _06751_ = sel_oi_one_hot_i[46] & i[239];
  assign _06762_ = i[255] & sel_oi_one_hot_i[47];
  assign _06772_ = _06762_ | _06751_;
  assign _06783_ = _06772_ | _06740_;
  assign _06794_ = _06783_ | _06708_;
  assign o[47] = _06794_ | _06633_;
  assign _06814_ = sel_oi_one_hot_i[32] & i[14];
  assign _06825_ = sel_oi_one_hot_i[33] & i[30];
  assign _06835_ = _06825_ | _06814_;
  assign _06846_ = sel_oi_one_hot_i[34] & i[46];
  assign _06857_ = sel_oi_one_hot_i[35] & i[62];
  assign _06867_ = _06857_ | _06846_;
  assign _06878_ = _06867_ | _06835_;
  assign _06889_ = sel_oi_one_hot_i[36] & i[78];
  assign _06899_ = sel_oi_one_hot_i[37] & i[94];
  assign _06910_ = _06899_ | _06889_;
  assign _06921_ = sel_oi_one_hot_i[38] & i[110];
  assign _06931_ = sel_oi_one_hot_i[39] & i[126];
  assign _06942_ = _06931_ | _06921_;
  assign _06953_ = _06942_ | _06910_;
  assign _06963_ = _06953_ | _06878_;
  assign _06974_ = sel_oi_one_hot_i[40] & i[142];
  assign _06985_ = sel_oi_one_hot_i[41] & i[158];
  assign _06995_ = _06985_ | _06974_;
  assign _07006_ = sel_oi_one_hot_i[42] & i[174];
  assign _07017_ = sel_oi_one_hot_i[43] & i[190];
  assign _07027_ = _07017_ | _07006_;
  assign _07038_ = _07027_ | _06995_;
  assign _07049_ = sel_oi_one_hot_i[44] & i[206];
  assign _07059_ = sel_oi_one_hot_i[45] & i[222];
  assign _07070_ = _07059_ | _07049_;
  assign _07081_ = sel_oi_one_hot_i[46] & i[238];
  assign _07092_ = i[254] & sel_oi_one_hot_i[47];
  assign _07102_ = _07092_ | _07081_;
  assign _07113_ = _07102_ | _07070_;
  assign _07124_ = _07113_ | _07038_;
  assign o[46] = _07124_ | _06963_;
  assign _07144_ = sel_oi_one_hot_i[0] & i[15];
  assign _07155_ = sel_oi_one_hot_i[1] & i[31];
  assign _07165_ = _07155_ | _07144_;
  assign _07176_ = sel_oi_one_hot_i[2] & i[47];
  assign _07187_ = sel_oi_one_hot_i[3] & i[63];
  assign _07197_ = _07187_ | _07176_;
  assign _07208_ = _07197_ | _07165_;
  assign _07219_ = sel_oi_one_hot_i[4] & i[79];
  assign _07229_ = sel_oi_one_hot_i[5] & i[95];
  assign _07240_ = _07229_ | _07219_;
  assign _07251_ = sel_oi_one_hot_i[6] & i[111];
  assign _07261_ = sel_oi_one_hot_i[7] & i[127];
  assign _07272_ = _07261_ | _07251_;
  assign _07283_ = _07272_ | _07240_;
  assign _07293_ = _07283_ | _07208_;
  assign _07304_ = sel_oi_one_hot_i[8] & i[143];
  assign _07315_ = sel_oi_one_hot_i[9] & i[159];
  assign _07325_ = _07315_ | _07304_;
  assign _07336_ = sel_oi_one_hot_i[10] & i[175];
  assign _07347_ = sel_oi_one_hot_i[11] & i[191];
  assign _07357_ = _07347_ | _07336_;
  assign _07368_ = _07357_ | _07325_;
  assign _07379_ = sel_oi_one_hot_i[12] & i[207];
  assign _07389_ = sel_oi_one_hot_i[13] & i[223];
  assign _07400_ = _07389_ | _07379_;
  assign _07411_ = sel_oi_one_hot_i[14] & i[239];
  assign _07422_ = sel_oi_one_hot_i[15] & i[255];
  assign _07432_ = _07422_ | _07411_;
  assign _07443_ = _07432_ | _07400_;
  assign _07454_ = _07443_ | _07368_;
  assign o[15] = _07454_ | _07293_;
  assign _07474_ = sel_oi_one_hot_i[32] & i[13];
  assign _07485_ = sel_oi_one_hot_i[33] & i[29];
  assign _07495_ = _07485_ | _07474_;
  assign _07506_ = sel_oi_one_hot_i[34] & i[45];
  assign _07517_ = sel_oi_one_hot_i[35] & i[61];
  assign _07527_ = _07517_ | _07506_;
  assign _07538_ = _07527_ | _07495_;
  assign _07549_ = sel_oi_one_hot_i[36] & i[77];
  assign _07554_ = sel_oi_one_hot_i[37] & i[93];
  assign _07555_ = _07554_ | _07549_;
  assign _07556_ = sel_oi_one_hot_i[38] & i[109];
  assign _07557_ = sel_oi_one_hot_i[39] & i[125];
  assign _07558_ = _07557_ | _07556_;
  assign _07559_ = _07558_ | _07555_;
  assign _07560_ = _07559_ | _07538_;
  assign _07561_ = sel_oi_one_hot_i[40] & i[141];
  assign _07562_ = sel_oi_one_hot_i[41] & i[157];
  assign _07563_ = _07562_ | _07561_;
  assign _07564_ = sel_oi_one_hot_i[42] & i[173];
  assign _07565_ = sel_oi_one_hot_i[43] & i[189];
  assign _07566_ = _07565_ | _07564_;
  assign _07567_ = _07566_ | _07563_;
  assign _07568_ = sel_oi_one_hot_i[44] & i[205];
  assign _07569_ = sel_oi_one_hot_i[45] & i[221];
  assign _07570_ = _07569_ | _07568_;
  assign _07571_ = sel_oi_one_hot_i[46] & i[237];
  assign _07572_ = i[253] & sel_oi_one_hot_i[47];
  assign _07573_ = _07572_ | _07571_;
  assign _07574_ = _07573_ | _07570_;
  assign _07575_ = _07574_ | _07567_;
  assign o[45] = _07575_ | _07560_;
  assign _07576_ = sel_oi_one_hot_i[32] & i[12];
  assign _07577_ = sel_oi_one_hot_i[33] & i[28];
  assign _07578_ = _07577_ | _07576_;
  assign _07579_ = sel_oi_one_hot_i[34] & i[44];
  assign _07580_ = sel_oi_one_hot_i[35] & i[60];
  assign _07581_ = _07580_ | _07579_;
  assign _07582_ = _07581_ | _07578_;
  assign _07583_ = sel_oi_one_hot_i[36] & i[76];
  assign _07584_ = sel_oi_one_hot_i[37] & i[92];
  assign _07585_ = _07584_ | _07583_;
  assign _07586_ = sel_oi_one_hot_i[38] & i[108];
  assign _07587_ = sel_oi_one_hot_i[39] & i[124];
  assign _07588_ = _07587_ | _07586_;
  assign _07589_ = _07588_ | _07585_;
  assign _07590_ = _07589_ | _07582_;
  assign _07591_ = sel_oi_one_hot_i[40] & i[140];
  assign _07592_ = sel_oi_one_hot_i[41] & i[156];
  assign _07593_ = _07592_ | _07591_;
  assign _07594_ = sel_oi_one_hot_i[42] & i[172];
  assign _07595_ = sel_oi_one_hot_i[43] & i[188];
  assign _07596_ = _07595_ | _07594_;
  assign _07597_ = _07596_ | _07593_;
  assign _07598_ = sel_oi_one_hot_i[44] & i[204];
  assign _07599_ = sel_oi_one_hot_i[45] & i[220];
  assign _07600_ = _07599_ | _07598_;
  assign _07601_ = sel_oi_one_hot_i[46] & i[236];
  assign _07602_ = i[252] & sel_oi_one_hot_i[47];
  assign _07603_ = _07602_ | _07601_;
  assign _07604_ = _07603_ | _07600_;
  assign _07605_ = _07604_ | _07597_;
  assign o[44] = _07605_ | _07590_;
  assign _07606_ = sel_oi_one_hot_i[32] & i[11];
  assign _07607_ = sel_oi_one_hot_i[33] & i[27];
  assign _07608_ = _07607_ | _07606_;
  assign _07609_ = sel_oi_one_hot_i[34] & i[43];
  assign _07610_ = sel_oi_one_hot_i[35] & i[59];
  assign _07611_ = _07610_ | _07609_;
  assign _07612_ = _07611_ | _07608_;
  assign _07613_ = sel_oi_one_hot_i[36] & i[75];
  assign _07614_ = sel_oi_one_hot_i[37] & i[91];
  assign _07615_ = _07614_ | _07613_;
  assign _07616_ = sel_oi_one_hot_i[38] & i[107];
  assign _07617_ = sel_oi_one_hot_i[39] & i[123];
  assign _07618_ = _07617_ | _07616_;
  assign _07619_ = _07618_ | _07615_;
  assign _07620_ = _07619_ | _07612_;
  assign _07621_ = sel_oi_one_hot_i[40] & i[139];
  assign _07622_ = sel_oi_one_hot_i[41] & i[155];
  assign _07623_ = _07622_ | _07621_;
  assign _07624_ = sel_oi_one_hot_i[42] & i[171];
  assign _07625_ = sel_oi_one_hot_i[43] & i[187];
  assign _07626_ = _07625_ | _07624_;
  assign _07627_ = _07626_ | _07623_;
  assign _07628_ = sel_oi_one_hot_i[44] & i[203];
  assign _07629_ = sel_oi_one_hot_i[45] & i[219];
  assign _07630_ = _07629_ | _07628_;
  assign _07631_ = sel_oi_one_hot_i[46] & i[235];
  assign _07632_ = i[251] & sel_oi_one_hot_i[47];
  assign _07633_ = _07632_ | _07631_;
  assign _07634_ = _07633_ | _07630_;
  assign _07635_ = _07634_ | _07627_;
  assign o[43] = _07635_ | _07620_;
  assign _07636_ = sel_oi_one_hot_i[32] & i[10];
  assign _07637_ = sel_oi_one_hot_i[33] & i[26];
  assign _07638_ = _07637_ | _07636_;
  assign _07639_ = sel_oi_one_hot_i[34] & i[42];
  assign _07640_ = sel_oi_one_hot_i[35] & i[58];
  assign _07641_ = _07640_ | _07639_;
  assign _07642_ = _07641_ | _07638_;
  assign _07643_ = sel_oi_one_hot_i[36] & i[74];
  assign _07644_ = sel_oi_one_hot_i[37] & i[90];
  assign _07645_ = _07644_ | _07643_;
  assign _07646_ = sel_oi_one_hot_i[38] & i[106];
  assign _07647_ = sel_oi_one_hot_i[39] & i[122];
  assign _07648_ = _07647_ | _07646_;
  assign _07649_ = _07648_ | _07645_;
  assign _07650_ = _07649_ | _07642_;
  assign _07651_ = sel_oi_one_hot_i[40] & i[138];
  assign _07652_ = sel_oi_one_hot_i[41] & i[154];
  assign _07653_ = _07652_ | _07651_;
  assign _07654_ = sel_oi_one_hot_i[42] & i[170];
  assign _07655_ = sel_oi_one_hot_i[43] & i[186];
  assign _07656_ = _07655_ | _07654_;
  assign _07657_ = _07656_ | _07653_;
  assign _07658_ = sel_oi_one_hot_i[44] & i[202];
  assign _07659_ = sel_oi_one_hot_i[45] & i[218];
  assign _07660_ = _07659_ | _07658_;
  assign _07661_ = sel_oi_one_hot_i[46] & i[234];
  assign _07662_ = i[250] & sel_oi_one_hot_i[47];
  assign _07663_ = _07662_ | _07661_;
  assign _07664_ = _07663_ | _07660_;
  assign _07665_ = _07664_ | _07657_;
  assign o[42] = _07665_ | _07650_;
  assign _07666_ = sel_oi_one_hot_i[32] & i[9];
  assign _07667_ = sel_oi_one_hot_i[33] & i[25];
  assign _07668_ = _07667_ | _07666_;
  assign _07669_ = sel_oi_one_hot_i[34] & i[41];
  assign _07670_ = sel_oi_one_hot_i[35] & i[57];
  assign _07671_ = _07670_ | _07669_;
  assign _07672_ = _07671_ | _07668_;
  assign _07673_ = sel_oi_one_hot_i[36] & i[73];
  assign _07674_ = sel_oi_one_hot_i[37] & i[89];
  assign _07675_ = _07674_ | _07673_;
  assign _07676_ = sel_oi_one_hot_i[38] & i[105];
  assign _07677_ = sel_oi_one_hot_i[39] & i[121];
  assign _07678_ = _07677_ | _07676_;
  assign _07679_ = _07678_ | _07675_;
  assign _00000_ = _07679_ | _07672_;
  assign _00001_ = sel_oi_one_hot_i[40] & i[137];
  assign _00002_ = sel_oi_one_hot_i[41] & i[153];
  assign _00003_ = _00002_ | _00001_;
  assign _00004_ = sel_oi_one_hot_i[42] & i[169];
  assign _00005_ = sel_oi_one_hot_i[43] & i[185];
  assign _00006_ = _00005_ | _00004_;
  assign _00007_ = _00006_ | _00003_;
  assign _00008_ = sel_oi_one_hot_i[44] & i[201];
  assign _00009_ = sel_oi_one_hot_i[45] & i[217];
  assign _00010_ = _00009_ | _00008_;
  assign _00011_ = i[233] & sel_oi_one_hot_i[46];
  assign _00012_ = i[249] & sel_oi_one_hot_i[47];
  assign _00013_ = _00012_ | _00011_;
  assign _00014_ = _00013_ | _00010_;
  assign _00015_ = _00014_ | _00007_;
  assign o[41] = _00015_ | _00000_;
  assign _00016_ = sel_oi_one_hot_i[32] & i[8];
  assign _00017_ = sel_oi_one_hot_i[33] & i[24];
  assign _00018_ = _00017_ | _00016_;
  assign _00019_ = sel_oi_one_hot_i[34] & i[40];
  assign _00020_ = sel_oi_one_hot_i[35] & i[56];
  assign _00021_ = _00020_ | _00019_;
  assign _00022_ = _00021_ | _00018_;
  assign _00023_ = sel_oi_one_hot_i[36] & i[72];
  assign _00024_ = sel_oi_one_hot_i[37] & i[88];
  assign _00025_ = _00024_ | _00023_;
  assign _00026_ = sel_oi_one_hot_i[38] & i[104];
  assign _00027_ = sel_oi_one_hot_i[39] & i[120];
  assign _00028_ = _00027_ | _00026_;
  assign _00029_ = _00028_ | _00025_;
  assign _00030_ = _00029_ | _00022_;
  assign _00031_ = sel_oi_one_hot_i[40] & i[136];
  assign _00032_ = sel_oi_one_hot_i[41] & i[152];
  assign _00033_ = _00032_ | _00031_;
  assign _00034_ = sel_oi_one_hot_i[42] & i[168];
  assign _00035_ = sel_oi_one_hot_i[43] & i[184];
  assign _00036_ = _00035_ | _00034_;
  assign _00037_ = _00036_ | _00033_;
  assign _00038_ = sel_oi_one_hot_i[44] & i[200];
  assign _00039_ = sel_oi_one_hot_i[45] & i[216];
  assign _00040_ = _00039_ | _00038_;
  assign _00041_ = i[232] & sel_oi_one_hot_i[46];
  assign _00042_ = i[248] & sel_oi_one_hot_i[47];
  assign _00043_ = _00042_ | _00041_;
  assign _00044_ = _00043_ | _00040_;
  assign _00045_ = _00044_ | _00037_;
  assign o[40] = _00045_ | _00030_;
  assign _00046_ = sel_oi_one_hot_i[32] & i[7];
  assign _00047_ = sel_oi_one_hot_i[33] & i[23];
  assign _00048_ = _00047_ | _00046_;
  assign _00049_ = sel_oi_one_hot_i[34] & i[39];
  assign _00050_ = sel_oi_one_hot_i[35] & i[55];
  assign _00051_ = _00050_ | _00049_;
  assign _00052_ = _00051_ | _00048_;
  assign _00053_ = sel_oi_one_hot_i[36] & i[71];
  assign _00054_ = sel_oi_one_hot_i[37] & i[87];
  assign _00055_ = _00054_ | _00053_;
  assign _00056_ = sel_oi_one_hot_i[38] & i[103];
  assign _00057_ = sel_oi_one_hot_i[39] & i[119];
  assign _00058_ = _00057_ | _00056_;
  assign _00059_ = _00058_ | _00055_;
  assign _00060_ = _00059_ | _00052_;
  assign _00061_ = sel_oi_one_hot_i[40] & i[135];
  assign _00062_ = sel_oi_one_hot_i[41] & i[151];
  assign _00063_ = _00062_ | _00061_;
  assign _00064_ = sel_oi_one_hot_i[42] & i[167];
  assign _00065_ = sel_oi_one_hot_i[43] & i[183];
  assign _00066_ = _00065_ | _00064_;
  assign _00067_ = _00066_ | _00063_;
  assign _00068_ = sel_oi_one_hot_i[44] & i[199];
  assign _00069_ = sel_oi_one_hot_i[45] & i[215];
  assign _00070_ = _00069_ | _00068_;
  assign _00071_ = i[231] & sel_oi_one_hot_i[46];
  assign _00072_ = i[247] & sel_oi_one_hot_i[47];
  assign _00073_ = _00072_ | _00071_;
  assign _00074_ = _00073_ | _00070_;
  assign _00075_ = _00074_ | _00067_;
  assign o[39] = _00075_ | _00060_;
  assign _00076_ = sel_oi_one_hot_i[32] & i[6];
  assign _00077_ = sel_oi_one_hot_i[33] & i[22];
  assign _00078_ = _00077_ | _00076_;
  assign _00079_ = sel_oi_one_hot_i[34] & i[38];
  assign _00080_ = sel_oi_one_hot_i[35] & i[54];
  assign _00081_ = _00080_ | _00079_;
  assign _00082_ = _00081_ | _00078_;
  assign _00083_ = sel_oi_one_hot_i[36] & i[70];
  assign _00084_ = sel_oi_one_hot_i[37] & i[86];
  assign _00085_ = _00084_ | _00083_;
  assign _00086_ = sel_oi_one_hot_i[38] & i[102];
  assign _00087_ = sel_oi_one_hot_i[39] & i[118];
  assign _00088_ = _00087_ | _00086_;
  assign _00089_ = _00088_ | _00085_;
  assign _00090_ = _00089_ | _00082_;
  assign _00091_ = sel_oi_one_hot_i[40] & i[134];
  assign _00092_ = sel_oi_one_hot_i[41] & i[150];
  assign _00093_ = _00092_ | _00091_;
  assign _00094_ = sel_oi_one_hot_i[42] & i[166];
  assign _00095_ = sel_oi_one_hot_i[43] & i[182];
  assign _00096_ = _00095_ | _00094_;
  assign _00097_ = _00096_ | _00093_;
  assign _00098_ = sel_oi_one_hot_i[44] & i[198];
  assign _00099_ = sel_oi_one_hot_i[45] & i[214];
  assign _00100_ = _00099_ | _00098_;
  assign _00101_ = i[230] & sel_oi_one_hot_i[46];
  assign _00102_ = i[246] & sel_oi_one_hot_i[47];
  assign _00103_ = _00102_ | _00101_;
  assign _00104_ = _00103_ | _00100_;
  assign _00105_ = _00104_ | _00097_;
  assign o[38] = _00105_ | _00090_;
  assign _00106_ = sel_oi_one_hot_i[32] & i[5];
  assign _00107_ = sel_oi_one_hot_i[33] & i[21];
  assign _00108_ = _00107_ | _00106_;
  assign _00109_ = sel_oi_one_hot_i[34] & i[37];
  assign _00110_ = sel_oi_one_hot_i[35] & i[53];
  assign _00111_ = _00110_ | _00109_;
  assign _00112_ = _00111_ | _00108_;
  assign _00113_ = sel_oi_one_hot_i[36] & i[69];
  assign _00114_ = sel_oi_one_hot_i[37] & i[85];
  assign _00115_ = _00114_ | _00113_;
  assign _00116_ = sel_oi_one_hot_i[38] & i[101];
  assign _00117_ = sel_oi_one_hot_i[39] & i[117];
  assign _00118_ = _00117_ | _00116_;
  assign _00119_ = _00118_ | _00115_;
  assign _00120_ = _00119_ | _00112_;
  assign _00121_ = sel_oi_one_hot_i[40] & i[133];
  assign _00122_ = sel_oi_one_hot_i[41] & i[149];
  assign _00123_ = _00122_ | _00121_;
  assign _00124_ = sel_oi_one_hot_i[42] & i[165];
  assign _00125_ = sel_oi_one_hot_i[43] & i[181];
  assign _00126_ = _00125_ | _00124_;
  assign _00127_ = _00126_ | _00123_;
  assign _00128_ = sel_oi_one_hot_i[44] & i[197];
  assign _00129_ = sel_oi_one_hot_i[45] & i[213];
  assign _00130_ = _00129_ | _00128_;
  assign _00131_ = i[229] & sel_oi_one_hot_i[46];
  assign _00132_ = i[245] & sel_oi_one_hot_i[47];
  assign _00133_ = _00132_ | _00131_;
  assign _00134_ = _00133_ | _00130_;
  assign _00135_ = _00134_ | _00127_;
  assign o[37] = _00135_ | _00120_;
  assign _00136_ = sel_oi_one_hot_i[32] & i[4];
  assign _00137_ = sel_oi_one_hot_i[33] & i[20];
  assign _00138_ = _00137_ | _00136_;
  assign _00139_ = sel_oi_one_hot_i[34] & i[36];
  assign _00140_ = sel_oi_one_hot_i[35] & i[52];
  assign _00141_ = _00140_ | _00139_;
  assign _00142_ = _00141_ | _00138_;
  assign _00143_ = sel_oi_one_hot_i[36] & i[68];
  assign _00144_ = sel_oi_one_hot_i[37] & i[84];
  assign _00145_ = _00144_ | _00143_;
  assign _00146_ = sel_oi_one_hot_i[38] & i[100];
  assign _00147_ = sel_oi_one_hot_i[39] & i[116];
  assign _00148_ = _00147_ | _00146_;
  assign _00149_ = _00148_ | _00145_;
  assign _00150_ = _00149_ | _00142_;
  assign _00151_ = sel_oi_one_hot_i[40] & i[132];
  assign _00152_ = sel_oi_one_hot_i[41] & i[148];
  assign _00153_ = _00152_ | _00151_;
  assign _00154_ = sel_oi_one_hot_i[42] & i[164];
  assign _00155_ = sel_oi_one_hot_i[43] & i[180];
  assign _00156_ = _00155_ | _00154_;
  assign _00157_ = _00156_ | _00153_;
  assign _00158_ = sel_oi_one_hot_i[44] & i[196];
  assign _00159_ = sel_oi_one_hot_i[45] & i[212];
  assign _00160_ = _00159_ | _00158_;
  assign _00161_ = i[228] & sel_oi_one_hot_i[46];
  assign _00162_ = i[244] & sel_oi_one_hot_i[47];
  assign _00163_ = _00162_ | _00161_;
  assign _00164_ = _00163_ | _00160_;
  assign _00165_ = _00164_ | _00157_;
  assign o[36] = _00165_ | _00150_;
  assign _00166_ = sel_oi_one_hot_i[0] & i[14];
  assign _00167_ = sel_oi_one_hot_i[1] & i[30];
  assign _00168_ = _00167_ | _00166_;
  assign _00169_ = sel_oi_one_hot_i[2] & i[46];
  assign _00170_ = sel_oi_one_hot_i[3] & i[62];
  assign _00171_ = _00170_ | _00169_;
  assign _00172_ = _00171_ | _00168_;
  assign _00173_ = sel_oi_one_hot_i[4] & i[78];
  assign _00174_ = sel_oi_one_hot_i[5] & i[94];
  assign _00175_ = _00174_ | _00173_;
  assign _00176_ = sel_oi_one_hot_i[6] & i[110];
  assign _00177_ = sel_oi_one_hot_i[7] & i[126];
  assign _00178_ = _00177_ | _00176_;
  assign _00179_ = _00178_ | _00175_;
  assign _00180_ = _00179_ | _00172_;
  assign _00181_ = sel_oi_one_hot_i[8] & i[142];
  assign _00182_ = sel_oi_one_hot_i[9] & i[158];
  assign _00183_ = _00182_ | _00181_;
  assign _00184_ = sel_oi_one_hot_i[10] & i[174];
  assign _00185_ = sel_oi_one_hot_i[11] & i[190];
  assign _00186_ = _00185_ | _00184_;
  assign _00187_ = _00186_ | _00183_;
  assign _00188_ = sel_oi_one_hot_i[12] & i[206];
  assign _00189_ = sel_oi_one_hot_i[13] & i[222];
  assign _00190_ = _00189_ | _00188_;
  assign _00191_ = sel_oi_one_hot_i[14] & i[238];
  assign _00192_ = sel_oi_one_hot_i[15] & i[254];
  assign _00193_ = _00192_ | _00191_;
  assign _00194_ = _00193_ | _00190_;
  assign _00195_ = _00194_ | _00187_;
  assign o[14] = _00195_ | _00180_;
  assign _00196_ = sel_oi_one_hot_i[32] & i[3];
  assign _00197_ = sel_oi_one_hot_i[33] & i[19];
  assign _00198_ = _00197_ | _00196_;
  assign _00199_ = sel_oi_one_hot_i[34] & i[35];
  assign _00200_ = sel_oi_one_hot_i[35] & i[51];
  assign _00201_ = _00200_ | _00199_;
  assign _00202_ = _00201_ | _00198_;
  assign _00203_ = sel_oi_one_hot_i[36] & i[67];
  assign _00204_ = sel_oi_one_hot_i[37] & i[83];
  assign _00205_ = _00204_ | _00203_;
  assign _00206_ = sel_oi_one_hot_i[38] & i[99];
  assign _00207_ = sel_oi_one_hot_i[39] & i[115];
  assign _00208_ = _00207_ | _00206_;
  assign _00209_ = _00208_ | _00205_;
  assign _00210_ = _00209_ | _00202_;
  assign _00211_ = sel_oi_one_hot_i[40] & i[131];
  assign _00212_ = sel_oi_one_hot_i[41] & i[147];
  assign _00213_ = _00212_ | _00211_;
  assign _00214_ = sel_oi_one_hot_i[42] & i[163];
  assign _00215_ = sel_oi_one_hot_i[43] & i[179];
  assign _00216_ = _00215_ | _00214_;
  assign _00217_ = _00216_ | _00213_;
  assign _00218_ = sel_oi_one_hot_i[44] & i[195];
  assign _00219_ = sel_oi_one_hot_i[45] & i[211];
  assign _00220_ = _00219_ | _00218_;
  assign _00221_ = i[227] & sel_oi_one_hot_i[46];
  assign _00222_ = i[243] & sel_oi_one_hot_i[47];
  assign _00223_ = _00222_ | _00221_;
  assign _00224_ = _00223_ | _00220_;
  assign _00225_ = _00224_ | _00217_;
  assign o[35] = _00225_ | _00210_;
  assign _00226_ = sel_oi_one_hot_i[32] & i[2];
  assign _00227_ = sel_oi_one_hot_i[33] & i[18];
  assign _00228_ = _00227_ | _00226_;
  assign _00229_ = sel_oi_one_hot_i[34] & i[34];
  assign _00230_ = sel_oi_one_hot_i[35] & i[50];
  assign _00231_ = _00230_ | _00229_;
  assign _00232_ = _00231_ | _00228_;
  assign _00233_ = sel_oi_one_hot_i[36] & i[66];
  assign _00234_ = sel_oi_one_hot_i[37] & i[82];
  assign _00235_ = _00234_ | _00233_;
  assign _00236_ = sel_oi_one_hot_i[38] & i[98];
  assign _00237_ = sel_oi_one_hot_i[39] & i[114];
  assign _00238_ = _00237_ | _00236_;
  assign _00239_ = _00238_ | _00235_;
  assign _00240_ = _00239_ | _00232_;
  assign _00241_ = sel_oi_one_hot_i[40] & i[130];
  assign _00242_ = sel_oi_one_hot_i[41] & i[146];
  assign _00243_ = _00242_ | _00241_;
  assign _00244_ = sel_oi_one_hot_i[42] & i[162];
  assign _00245_ = sel_oi_one_hot_i[43] & i[178];
  assign _00246_ = _00245_ | _00244_;
  assign _00247_ = _00246_ | _00243_;
  assign _00248_ = sel_oi_one_hot_i[44] & i[194];
  assign _00249_ = sel_oi_one_hot_i[45] & i[210];
  assign _00250_ = _00249_ | _00248_;
  assign _00251_ = i[226] & sel_oi_one_hot_i[46];
  assign _00252_ = i[242] & sel_oi_one_hot_i[47];
  assign _00253_ = _00252_ | _00251_;
  assign _00254_ = _00253_ | _00250_;
  assign _00255_ = _00254_ | _00247_;
  assign o[34] = _00255_ | _00240_;
  assign _00256_ = sel_oi_one_hot_i[32] & i[1];
  assign _00257_ = sel_oi_one_hot_i[33] & i[17];
  assign _00258_ = _00257_ | _00256_;
  assign _00259_ = sel_oi_one_hot_i[34] & i[33];
  assign _00260_ = sel_oi_one_hot_i[35] & i[49];
  assign _00261_ = _00260_ | _00259_;
  assign _00262_ = _00261_ | _00258_;
  assign _00263_ = sel_oi_one_hot_i[36] & i[65];
  assign _00264_ = sel_oi_one_hot_i[37] & i[81];
  assign _00265_ = _00264_ | _00263_;
  assign _00266_ = sel_oi_one_hot_i[38] & i[97];
  assign _00267_ = sel_oi_one_hot_i[39] & i[113];
  assign _00268_ = _00267_ | _00266_;
  assign _00269_ = _00268_ | _00265_;
  assign _00270_ = _00269_ | _00262_;
  assign _00271_ = sel_oi_one_hot_i[40] & i[129];
  assign _00272_ = sel_oi_one_hot_i[41] & i[145];
  assign _00273_ = _00272_ | _00271_;
  assign _00274_ = sel_oi_one_hot_i[42] & i[161];
  assign _00275_ = sel_oi_one_hot_i[43] & i[177];
  assign _00276_ = _00275_ | _00274_;
  assign _00277_ = _00276_ | _00273_;
  assign _00278_ = sel_oi_one_hot_i[44] & i[193];
  assign _00279_ = sel_oi_one_hot_i[45] & i[209];
  assign _00280_ = _00279_ | _00278_;
  assign _00281_ = i[225] & sel_oi_one_hot_i[46];
  assign _00282_ = i[241] & sel_oi_one_hot_i[47];
  assign _00283_ = _00282_ | _00281_;
  assign _00284_ = _00283_ | _00280_;
  assign _00285_ = _00284_ | _00277_;
  assign o[33] = _00285_ | _00270_;
  assign _00286_ = sel_oi_one_hot_i[32] & i[0];
  assign _00287_ = sel_oi_one_hot_i[33] & i[16];
  assign _00288_ = _00287_ | _00286_;
  assign _00289_ = sel_oi_one_hot_i[34] & i[32];
  assign _00290_ = sel_oi_one_hot_i[35] & i[48];
  assign _00291_ = _00290_ | _00289_;
  assign _00292_ = _00291_ | _00288_;
  assign _00293_ = sel_oi_one_hot_i[36] & i[64];
  assign _00294_ = sel_oi_one_hot_i[37] & i[80];
  assign _00295_ = _00294_ | _00293_;
  assign _00296_ = sel_oi_one_hot_i[38] & i[96];
  assign _00297_ = sel_oi_one_hot_i[39] & i[112];
  assign _00298_ = _00297_ | _00296_;
  assign _00299_ = _00298_ | _00295_;
  assign _00300_ = _00299_ | _00292_;
  assign _00301_ = sel_oi_one_hot_i[40] & i[128];
  assign _00302_ = sel_oi_one_hot_i[41] & i[144];
  assign _00303_ = _00302_ | _00301_;
  assign _00304_ = sel_oi_one_hot_i[42] & i[160];
  assign _00305_ = sel_oi_one_hot_i[43] & i[176];
  assign _00306_ = _00305_ | _00304_;
  assign _00307_ = _00306_ | _00303_;
  assign _00308_ = sel_oi_one_hot_i[44] & i[192];
  assign _00309_ = sel_oi_one_hot_i[45] & i[208];
  assign _00310_ = _00309_ | _00308_;
  assign _00311_ = sel_oi_one_hot_i[46] & i[224];
  assign _00312_ = sel_oi_one_hot_i[47] & i[240];
  assign _00313_ = _00312_ | _00311_;
  assign _00314_ = _00313_ | _00310_;
  assign _00315_ = _00314_ | _00307_;
  assign o[32] = _00315_ | _00300_;
  assign _00316_ = sel_oi_one_hot_i[0] & i[13];
  assign _00317_ = sel_oi_one_hot_i[1] & i[29];
  assign _00318_ = _00317_ | _00316_;
  assign _00319_ = sel_oi_one_hot_i[2] & i[45];
  assign _00320_ = sel_oi_one_hot_i[3] & i[61];
  assign _00321_ = _00320_ | _00319_;
  assign _00322_ = _00321_ | _00318_;
  assign _00323_ = sel_oi_one_hot_i[4] & i[77];
  assign _00324_ = sel_oi_one_hot_i[5] & i[93];
  assign _00325_ = _00324_ | _00323_;
  assign _00326_ = sel_oi_one_hot_i[6] & i[109];
  assign _00327_ = sel_oi_one_hot_i[7] & i[125];
  assign _00328_ = _00327_ | _00326_;
  assign _00329_ = _00328_ | _00325_;
  assign _00330_ = _00329_ | _00322_;
  assign _00331_ = sel_oi_one_hot_i[8] & i[141];
  assign _00332_ = sel_oi_one_hot_i[9] & i[157];
  assign _00333_ = _00332_ | _00331_;
  assign _00334_ = sel_oi_one_hot_i[10] & i[173];
  assign _00335_ = sel_oi_one_hot_i[11] & i[189];
  assign _00336_ = _00335_ | _00334_;
  assign _00337_ = _00336_ | _00333_;
  assign _00338_ = sel_oi_one_hot_i[12] & i[205];
  assign _00339_ = sel_oi_one_hot_i[13] & i[221];
  assign _00340_ = _00339_ | _00338_;
  assign _00341_ = sel_oi_one_hot_i[14] & i[237];
  assign _00342_ = sel_oi_one_hot_i[15] & i[253];
  assign _00343_ = _00342_ | _00341_;
  assign _00344_ = _00343_ | _00340_;
  assign _00345_ = _00344_ | _00337_;
  assign o[13] = _00345_ | _00330_;
  assign _00346_ = sel_oi_one_hot_i[48] & i[15];
  assign _00347_ = sel_oi_one_hot_i[49] & i[31];
  assign _00348_ = _00347_ | _00346_;
  assign _00349_ = sel_oi_one_hot_i[50] & i[47];
  assign _00350_ = sel_oi_one_hot_i[51] & i[63];
  assign _00351_ = _00350_ | _00349_;
  assign _00352_ = _00351_ | _00348_;
  assign _00353_ = sel_oi_one_hot_i[52] & i[79];
  assign _00354_ = sel_oi_one_hot_i[53] & i[95];
  assign _00355_ = _00354_ | _00353_;
  assign _00356_ = sel_oi_one_hot_i[54] & i[111];
  assign _00357_ = sel_oi_one_hot_i[55] & i[127];
  assign _00358_ = _00357_ | _00356_;
  assign _00359_ = _00358_ | _00355_;
  assign _00360_ = _00359_ | _00352_;
  assign _00361_ = sel_oi_one_hot_i[56] & i[143];
  assign _00362_ = sel_oi_one_hot_i[57] & i[159];
  assign _00363_ = _00362_ | _00361_;
  assign _00364_ = sel_oi_one_hot_i[58] & i[175];
  assign _00365_ = sel_oi_one_hot_i[59] & i[191];
  assign _00366_ = _00365_ | _00364_;
  assign _00367_ = _00366_ | _00363_;
  assign _00368_ = sel_oi_one_hot_i[60] & i[207];
  assign _00369_ = sel_oi_one_hot_i[61] & i[223];
  assign _00370_ = _00369_ | _00368_;
  assign _00371_ = sel_oi_one_hot_i[62] & i[239];
  assign _00372_ = sel_oi_one_hot_i[63] & i[255];
  assign _00373_ = _00372_ | _00371_;
  assign _00374_ = _00373_ | _00370_;
  assign _00375_ = _00374_ | _00367_;
  assign o[63] = _00375_ | _00360_;
  assign _00376_ = sel_oi_one_hot_i[48] & i[14];
  assign _00377_ = sel_oi_one_hot_i[49] & i[30];
  assign _00378_ = _00377_ | _00376_;
  assign _00379_ = sel_oi_one_hot_i[50] & i[46];
  assign _00380_ = sel_oi_one_hot_i[51] & i[62];
  assign _00381_ = _00380_ | _00379_;
  assign _00382_ = _00381_ | _00378_;
  assign _00383_ = sel_oi_one_hot_i[52] & i[78];
  assign _00384_ = sel_oi_one_hot_i[53] & i[94];
  assign _00385_ = _00384_ | _00383_;
  assign _00386_ = sel_oi_one_hot_i[54] & i[110];
  assign _00387_ = sel_oi_one_hot_i[55] & i[126];
  assign _00388_ = _00387_ | _00386_;
  assign _00389_ = _00388_ | _00385_;
  assign _00390_ = _00389_ | _00382_;
  assign _00391_ = sel_oi_one_hot_i[56] & i[142];
  assign _00392_ = sel_oi_one_hot_i[57] & i[158];
  assign _00393_ = _00392_ | _00391_;
  assign _00394_ = sel_oi_one_hot_i[58] & i[174];
  assign _00395_ = sel_oi_one_hot_i[59] & i[190];
  assign _00396_ = _00395_ | _00394_;
  assign _00397_ = _00396_ | _00393_;
  assign _00398_ = sel_oi_one_hot_i[60] & i[206];
  assign _00399_ = sel_oi_one_hot_i[61] & i[222];
  assign _00400_ = _00399_ | _00398_;
  assign _00401_ = sel_oi_one_hot_i[62] & i[238];
  assign _00402_ = sel_oi_one_hot_i[63] & i[254];
  assign _00403_ = _00402_ | _00401_;
  assign _00404_ = _00403_ | _00400_;
  assign _00405_ = _00404_ | _00397_;
  assign o[62] = _00405_ | _00390_;
  assign _00406_ = sel_oi_one_hot_i[48] & i[13];
  assign _00407_ = sel_oi_one_hot_i[49] & i[29];
  assign _00408_ = _00407_ | _00406_;
  assign _00409_ = sel_oi_one_hot_i[50] & i[45];
  assign _00410_ = sel_oi_one_hot_i[51] & i[61];
  assign _00411_ = _00410_ | _00409_;
  assign _00412_ = _00411_ | _00408_;
  assign _00413_ = sel_oi_one_hot_i[52] & i[77];
  assign _00414_ = sel_oi_one_hot_i[53] & i[93];
  assign _00415_ = _00414_ | _00413_;
  assign _00416_ = sel_oi_one_hot_i[54] & i[109];
  assign _00417_ = sel_oi_one_hot_i[55] & i[125];
  assign _00418_ = _00417_ | _00416_;
  assign _00419_ = _00418_ | _00415_;
  assign _00420_ = _00419_ | _00412_;
  assign _00421_ = sel_oi_one_hot_i[56] & i[141];
  assign _00422_ = sel_oi_one_hot_i[57] & i[157];
  assign _00423_ = _00422_ | _00421_;
  assign _00424_ = sel_oi_one_hot_i[58] & i[173];
  assign _00425_ = sel_oi_one_hot_i[59] & i[189];
  assign _00426_ = _00425_ | _00424_;
  assign _00427_ = _00426_ | _00423_;
  assign _00428_ = sel_oi_one_hot_i[60] & i[205];
  assign _00429_ = sel_oi_one_hot_i[61] & i[221];
  assign _00430_ = _00429_ | _00428_;
  assign _00431_ = sel_oi_one_hot_i[62] & i[237];
  assign _00432_ = sel_oi_one_hot_i[63] & i[253];
  assign _00433_ = _00432_ | _00431_;
  assign _00434_ = _00433_ | _00430_;
  assign _00435_ = _00434_ | _00427_;
  assign o[61] = _00435_ | _00420_;
  assign _00436_ = sel_oi_one_hot_i[0] & i[12];
  assign _00437_ = sel_oi_one_hot_i[1] & i[28];
  assign _00438_ = _00437_ | _00436_;
  assign _00439_ = sel_oi_one_hot_i[2] & i[44];
  assign _00440_ = sel_oi_one_hot_i[3] & i[60];
  assign _00441_ = _00440_ | _00439_;
  assign _00442_ = _00441_ | _00438_;
  assign _00443_ = sel_oi_one_hot_i[4] & i[76];
  assign _00444_ = sel_oi_one_hot_i[5] & i[92];
  assign _00445_ = _00444_ | _00443_;
  assign _00446_ = sel_oi_one_hot_i[6] & i[108];
  assign _00447_ = sel_oi_one_hot_i[7] & i[124];
  assign _00448_ = _00447_ | _00446_;
  assign _00449_ = _00448_ | _00445_;
  assign _00450_ = _00449_ | _00442_;
  assign _00451_ = sel_oi_one_hot_i[8] & i[140];
  assign _00452_ = sel_oi_one_hot_i[9] & i[156];
  assign _00453_ = _00452_ | _00451_;
  assign _00454_ = sel_oi_one_hot_i[10] & i[172];
  assign _00455_ = sel_oi_one_hot_i[11] & i[188];
  assign _00456_ = _00455_ | _00454_;
  assign _00457_ = _00456_ | _00453_;
  assign _00458_ = sel_oi_one_hot_i[12] & i[204];
  assign _00459_ = sel_oi_one_hot_i[13] & i[220];
  assign _00460_ = _00459_ | _00458_;
  assign _00461_ = sel_oi_one_hot_i[14] & i[236];
  assign _00462_ = sel_oi_one_hot_i[15] & i[252];
  assign _00463_ = _00462_ | _00461_;
  assign _00464_ = _00463_ | _00460_;
  assign _00465_ = _00464_ | _00457_;
  assign o[12] = _00465_ | _00450_;
  assign _00466_ = sel_oi_one_hot_i[48] & i[12];
  assign _00467_ = sel_oi_one_hot_i[49] & i[28];
  assign _00468_ = _00467_ | _00466_;
  assign _00469_ = sel_oi_one_hot_i[50] & i[44];
  assign _00470_ = sel_oi_one_hot_i[51] & i[60];
  assign _00471_ = _00470_ | _00469_;
  assign _00472_ = _00471_ | _00468_;
  assign _00473_ = sel_oi_one_hot_i[52] & i[76];
  assign _00474_ = sel_oi_one_hot_i[53] & i[92];
  assign _00475_ = _00474_ | _00473_;
  assign _00476_ = sel_oi_one_hot_i[54] & i[108];
  assign _00477_ = sel_oi_one_hot_i[55] & i[124];
  assign _00478_ = _00477_ | _00476_;
  assign _00479_ = _00478_ | _00475_;
  assign _00480_ = _00479_ | _00472_;
  assign _00481_ = sel_oi_one_hot_i[56] & i[140];
  assign _00482_ = sel_oi_one_hot_i[57] & i[156];
  assign _00483_ = _00482_ | _00481_;
  assign _00484_ = sel_oi_one_hot_i[58] & i[172];
  assign _00485_ = sel_oi_one_hot_i[59] & i[188];
  assign _00486_ = _00485_ | _00484_;
  assign _00487_ = _00486_ | _00483_;
  assign _00488_ = sel_oi_one_hot_i[60] & i[204];
  assign _00489_ = sel_oi_one_hot_i[61] & i[220];
  assign _00490_ = _00489_ | _00488_;
  assign _00491_ = sel_oi_one_hot_i[62] & i[236];
  assign _00492_ = sel_oi_one_hot_i[63] & i[252];
  assign _00493_ = _00492_ | _00491_;
  assign _00494_ = _00493_ | _00490_;
  assign _00495_ = _00494_ | _00487_;
  assign o[60] = _00495_ | _00480_;
  assign _00496_ = sel_oi_one_hot_i[48] & i[11];
  assign _00497_ = sel_oi_one_hot_i[49] & i[27];
  assign _00498_ = _00497_ | _00496_;
  assign _00499_ = sel_oi_one_hot_i[50] & i[43];
  assign _00500_ = sel_oi_one_hot_i[51] & i[59];
  assign _00501_ = _00500_ | _00499_;
  assign _00502_ = _00501_ | _00498_;
  assign _00503_ = sel_oi_one_hot_i[52] & i[75];
  assign _00504_ = sel_oi_one_hot_i[53] & i[91];
  assign _00505_ = _00504_ | _00503_;
  assign _00506_ = sel_oi_one_hot_i[54] & i[107];
  assign _00507_ = sel_oi_one_hot_i[55] & i[123];
  assign _00508_ = _00507_ | _00506_;
  assign _00509_ = _00508_ | _00505_;
  assign _00510_ = _00509_ | _00502_;
  assign _00511_ = sel_oi_one_hot_i[56] & i[139];
  assign _00512_ = sel_oi_one_hot_i[57] & i[155];
  assign _00513_ = _00512_ | _00511_;
  assign _00514_ = sel_oi_one_hot_i[58] & i[171];
  assign _00515_ = sel_oi_one_hot_i[59] & i[187];
  assign _00516_ = _00515_ | _00514_;
  assign _00517_ = _00516_ | _00513_;
  assign _00518_ = sel_oi_one_hot_i[60] & i[203];
  assign _00519_ = sel_oi_one_hot_i[61] & i[219];
  assign _00520_ = _00519_ | _00518_;
  assign _00521_ = sel_oi_one_hot_i[62] & i[235];
  assign _00522_ = sel_oi_one_hot_i[63] & i[251];
  assign _00523_ = _00522_ | _00521_;
  assign _00524_ = _00523_ | _00520_;
  assign _00525_ = _00524_ | _00517_;
  assign o[59] = _00525_ | _00510_;
  assign _00526_ = sel_oi_one_hot_i[48] & i[10];
  assign _00527_ = sel_oi_one_hot_i[49] & i[26];
  assign _00528_ = _00527_ | _00526_;
  assign _00529_ = sel_oi_one_hot_i[50] & i[42];
  assign _00530_ = sel_oi_one_hot_i[51] & i[58];
  assign _00531_ = _00530_ | _00529_;
  assign _00532_ = _00531_ | _00528_;
  assign _00533_ = sel_oi_one_hot_i[52] & i[74];
  assign _00534_ = sel_oi_one_hot_i[53] & i[90];
  assign _00535_ = _00534_ | _00533_;
  assign _00536_ = sel_oi_one_hot_i[54] & i[106];
  assign _00537_ = sel_oi_one_hot_i[55] & i[122];
  assign _00538_ = _00537_ | _00536_;
  assign _00539_ = _00538_ | _00535_;
  assign _00540_ = _00539_ | _00532_;
  assign _00541_ = sel_oi_one_hot_i[56] & i[138];
  assign _00542_ = sel_oi_one_hot_i[57] & i[154];
  assign _00543_ = _00542_ | _00541_;
  assign _00544_ = sel_oi_one_hot_i[58] & i[170];
  assign _00545_ = sel_oi_one_hot_i[59] & i[186];
  assign _00546_ = _00545_ | _00544_;
  assign _00547_ = _00546_ | _00543_;
  assign _00548_ = sel_oi_one_hot_i[60] & i[202];
  assign _00549_ = sel_oi_one_hot_i[61] & i[218];
  assign _00550_ = _00549_ | _00548_;
  assign _00551_ = sel_oi_one_hot_i[62] & i[234];
  assign _00552_ = sel_oi_one_hot_i[63] & i[250];
  assign _00553_ = _00552_ | _00551_;
  assign _00554_ = _00553_ | _00550_;
  assign _00555_ = _00554_ | _00547_;
  assign o[58] = _00555_ | _00540_;
  assign _00556_ = sel_oi_one_hot_i[48] & i[9];
  assign _00557_ = sel_oi_one_hot_i[49] & i[25];
  assign _00558_ = _00557_ | _00556_;
  assign _00559_ = sel_oi_one_hot_i[50] & i[41];
  assign _00560_ = sel_oi_one_hot_i[51] & i[57];
  assign _00561_ = _00560_ | _00559_;
  assign _00562_ = _00561_ | _00558_;
  assign _00563_ = sel_oi_one_hot_i[52] & i[73];
  assign _00564_ = sel_oi_one_hot_i[53] & i[89];
  assign _00565_ = _00564_ | _00563_;
  assign _00566_ = sel_oi_one_hot_i[54] & i[105];
  assign _00567_ = sel_oi_one_hot_i[55] & i[121];
  assign _00568_ = _00567_ | _00566_;
  assign _00569_ = _00568_ | _00565_;
  assign _00570_ = _00569_ | _00562_;
  assign _00571_ = sel_oi_one_hot_i[56] & i[137];
  assign _00572_ = sel_oi_one_hot_i[57] & i[153];
  assign _00573_ = _00572_ | _00571_;
  assign _00574_ = sel_oi_one_hot_i[58] & i[169];
  assign _00575_ = sel_oi_one_hot_i[59] & i[185];
  assign _00576_ = _00575_ | _00574_;
  assign _00577_ = _00576_ | _00573_;
  assign _00578_ = sel_oi_one_hot_i[60] & i[201];
  assign _00579_ = sel_oi_one_hot_i[61] & i[217];
  assign _00580_ = _00579_ | _00578_;
  assign _00581_ = sel_oi_one_hot_i[62] & i[233];
  assign _00582_ = sel_oi_one_hot_i[63] & i[249];
  assign _00583_ = _00582_ | _00581_;
  assign _00584_ = _00583_ | _00580_;
  assign _00585_ = _00584_ | _00577_;
  assign o[57] = _00585_ | _00570_;
  assign _00586_ = sel_oi_one_hot_i[48] & i[8];
  assign _00587_ = sel_oi_one_hot_i[49] & i[24];
  assign _00588_ = _00587_ | _00586_;
  assign _00589_ = sel_oi_one_hot_i[50] & i[40];
  assign _00590_ = sel_oi_one_hot_i[51] & i[56];
  assign _00591_ = _00590_ | _00589_;
  assign _00592_ = _00591_ | _00588_;
  assign _00593_ = sel_oi_one_hot_i[52] & i[72];
  assign _00594_ = sel_oi_one_hot_i[53] & i[88];
  assign _00595_ = _00594_ | _00593_;
  assign _00596_ = sel_oi_one_hot_i[54] & i[104];
  assign _00597_ = sel_oi_one_hot_i[55] & i[120];
  assign _00598_ = _00597_ | _00596_;
  assign _00599_ = _00598_ | _00595_;
  assign _00600_ = _00599_ | _00592_;
  assign _00601_ = sel_oi_one_hot_i[56] & i[136];
  assign _00602_ = sel_oi_one_hot_i[57] & i[152];
  assign _00603_ = _00602_ | _00601_;
  assign _00604_ = sel_oi_one_hot_i[58] & i[168];
  assign _00605_ = sel_oi_one_hot_i[59] & i[184];
  assign _00606_ = _00605_ | _00604_;
  assign _00607_ = _00606_ | _00603_;
  assign _00608_ = sel_oi_one_hot_i[60] & i[200];
  assign _00609_ = sel_oi_one_hot_i[61] & i[216];
  assign _00610_ = _00609_ | _00608_;
  assign _00611_ = sel_oi_one_hot_i[62] & i[232];
  assign _00612_ = sel_oi_one_hot_i[63] & i[248];
  assign _00613_ = _00612_ | _00611_;
  assign _00614_ = _00613_ | _00610_;
  assign _00615_ = _00614_ | _00607_;
  assign o[56] = _00615_ | _00600_;
  assign _00616_ = sel_oi_one_hot_i[48] & i[7];
  assign _00617_ = sel_oi_one_hot_i[49] & i[23];
  assign _00618_ = _00617_ | _00616_;
  assign _00619_ = sel_oi_one_hot_i[50] & i[39];
  assign _00620_ = sel_oi_one_hot_i[51] & i[55];
  assign _00621_ = _00620_ | _00619_;
  assign _00622_ = _00621_ | _00618_;
  assign _00623_ = sel_oi_one_hot_i[52] & i[71];
  assign _00624_ = sel_oi_one_hot_i[53] & i[87];
  assign _00625_ = _00624_ | _00623_;
  assign _00626_ = sel_oi_one_hot_i[54] & i[103];
  assign _00627_ = sel_oi_one_hot_i[55] & i[119];
  assign _00628_ = _00627_ | _00626_;
  assign _00629_ = _00628_ | _00625_;
  assign _00630_ = _00629_ | _00622_;
  assign _00631_ = sel_oi_one_hot_i[56] & i[135];
  assign _00632_ = sel_oi_one_hot_i[57] & i[151];
  assign _00633_ = _00632_ | _00631_;
  assign _00634_ = sel_oi_one_hot_i[58] & i[167];
  assign _00635_ = sel_oi_one_hot_i[59] & i[183];
  assign _00636_ = _00635_ | _00634_;
  assign _00637_ = _00636_ | _00633_;
  assign _00638_ = sel_oi_one_hot_i[60] & i[199];
  assign _00639_ = sel_oi_one_hot_i[61] & i[215];
  assign _00640_ = _00639_ | _00638_;
  assign _00641_ = sel_oi_one_hot_i[62] & i[231];
  assign _00642_ = sel_oi_one_hot_i[63] & i[247];
  assign _00643_ = _00642_ | _00641_;
  assign _00644_ = _00643_ | _00640_;
  assign _00645_ = _00644_ | _00637_;
  assign o[55] = _00645_ | _00630_;
  assign _00646_ = sel_oi_one_hot_i[48] & i[6];
  assign _00647_ = sel_oi_one_hot_i[49] & i[22];
  assign _00648_ = _00647_ | _00646_;
  assign _00649_ = sel_oi_one_hot_i[50] & i[38];
  assign _00650_ = sel_oi_one_hot_i[51] & i[54];
  assign _00651_ = _00650_ | _00649_;
  assign _00652_ = _00651_ | _00648_;
  assign _00653_ = sel_oi_one_hot_i[52] & i[70];
  assign _00654_ = sel_oi_one_hot_i[53] & i[86];
  assign _00655_ = _00654_ | _00653_;
  assign _00656_ = sel_oi_one_hot_i[54] & i[102];
  assign _00657_ = sel_oi_one_hot_i[55] & i[118];
  assign _00658_ = _00657_ | _00656_;
  assign _00659_ = _00658_ | _00655_;
  assign _00660_ = _00659_ | _00652_;
  assign _00661_ = sel_oi_one_hot_i[56] & i[134];
  assign _00662_ = sel_oi_one_hot_i[57] & i[150];
  assign _00663_ = _00662_ | _00661_;
  assign _00664_ = sel_oi_one_hot_i[58] & i[166];
  assign _00665_ = sel_oi_one_hot_i[59] & i[182];
  assign _00666_ = _00665_ | _00664_;
  assign _00667_ = _00666_ | _00663_;
  assign _00668_ = sel_oi_one_hot_i[60] & i[198];
  assign _00669_ = sel_oi_one_hot_i[61] & i[214];
  assign _00670_ = _00669_ | _00668_;
  assign _00671_ = sel_oi_one_hot_i[62] & i[230];
  assign _00672_ = sel_oi_one_hot_i[63] & i[246];
  assign _00673_ = _00672_ | _00671_;
  assign _00674_ = _00673_ | _00670_;
  assign _00675_ = _00674_ | _00667_;
  assign \l[0].mux_one_hot.data_i  = i;
  assign \l[0].mux_one_hot.data_o  = o[15:0];
  assign \l[0].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[15:0];
  assign \l[10].mux_one_hot.data_i  = i;
  assign \l[10].mux_one_hot.data_o  = o[175:160];
  assign \l[10].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[175:160];
  assign \l[11].mux_one_hot.data_i  = i;
  assign \l[11].mux_one_hot.data_o  = o[191:176];
  assign \l[11].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[191:176];
  assign \l[12].mux_one_hot.data_i  = i;
  assign \l[12].mux_one_hot.data_o  = o[207:192];
  assign \l[12].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[207:192];
  assign \l[13].mux_one_hot.data_i  = i;
  assign \l[13].mux_one_hot.data_o  = o[223:208];
  assign \l[13].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[223:208];
  assign \l[14].mux_one_hot.data_i  = i;
  assign \l[14].mux_one_hot.data_o  = o[239:224];
  assign \l[14].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[239:224];
  assign \l[15].mux_one_hot.data_i  = i;
  assign \l[15].mux_one_hot.data_o  = o[255:240];
  assign \l[15].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[255:240];
  assign \l[1].mux_one_hot.data_i  = i;
  assign \l[1].mux_one_hot.data_o  = o[31:16];
  assign \l[1].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[31:16];
  assign \l[2].mux_one_hot.data_i  = i;
  assign \l[2].mux_one_hot.data_o  = o[47:32];
  assign \l[2].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[47:32];
  assign \l[3].mux_one_hot.data_i  = i;
  assign \l[3].mux_one_hot.data_o  = o[63:48];
  assign \l[3].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[63:48];
  assign \l[4].mux_one_hot.data_i  = i;
  assign \l[4].mux_one_hot.data_o  = o[79:64];
  assign \l[4].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[79:64];
  assign \l[5].mux_one_hot.data_i  = i;
  assign \l[5].mux_one_hot.data_o  = o[95:80];
  assign \l[5].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[95:80];
  assign \l[6].mux_one_hot.data_i  = i;
  assign \l[6].mux_one_hot.data_o  = o[111:96];
  assign \l[6].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[111:96];
  assign \l[7].mux_one_hot.data_i  = i;
  assign \l[7].mux_one_hot.data_o  = o[127:112];
  assign \l[7].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[127:112];
  assign \l[8].mux_one_hot.data_i  = i;
  assign \l[8].mux_one_hot.data_o  = o[143:128];
  assign \l[8].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[143:128];
  assign \l[9].mux_one_hot.data_i  = i;
  assign \l[9].mux_one_hot.data_o  = o[159:144];
  assign \l[9].mux_one_hot.sel_one_hot_i  = sel_oi_one_hot_i[159:144];
endmodule
