module bsg_mux2_gatestack(i0, i1, i2, o);
  input [15:0] i0;
  wire [15:0] i0;
  input [15:0] i1;
  wire [15:0] i1;
  input [15:0] i2;
  wire [15:0] i2;
  output [15:0] o;
  wire [15:0] o;
  assign o[6] = i2[6] ? i1[6] : i0[6];
  assign o[7] = i2[7] ? i1[7] : i0[7];
  assign o[8] = i2[8] ? i1[8] : i0[8];
  assign o[9] = i2[9] ? i1[9] : i0[9];
  assign o[10] = i2[10] ? i1[10] : i0[10];
  assign o[11] = i2[11] ? i1[11] : i0[11];
  assign o[12] = i2[12] ? i1[12] : i0[12];
  assign o[13] = i2[13] ? i1[13] : i0[13];
  assign o[14] = i2[14] ? i1[14] : i0[14];
  assign o[15] = i2[15] ? i1[15] : i0[15];
  assign o[0] = i2[0] ? i1[0] : i0[0];
  assign o[1] = i2[1] ? i1[1] : i0[1];
  assign o[2] = i2[2] ? i1[2] : i0[2];
  assign o[3] = i2[3] ? i1[3] : i0[3];
  assign o[4] = i2[4] ? i1[4] : i0[4];
  assign o[5] = i2[5] ? i1[5] : i0[5];
endmodule
