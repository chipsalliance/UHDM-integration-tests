module bsg_counter_set_down(clk_i, reset_i, set_i, val_i, down_i, count_r_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  input clk_i;
  wire clk_i;
  output [15:0] count_r_o;
  wire [15:0] count_r_o;
  wire [15:0] ctr_n;
  reg [15:0] ctr_r;
  input down_i;
  wire down_i;
  input reset_i;
  wire reset_i;
  input set_i;
  wire set_i;
  input [15:0] val_i;
  wire [15:0] val_i;
  assign _033_ = set_i ? val_i[0] : ctr_r[0];
  assign ctr_n[0] = _033_ ^ down_i;
  assign _034_ = set_i ? val_i[1] : ctr_r[1];
  assign _035_ = ~(_034_ ^ _033_);
  assign ctr_n[1] = down_i ? _035_ : _034_;
  assign _036_ = set_i ? val_i[2] : ctr_r[2];
  assign _037_ = ~_036_;
  assign _038_ = _034_ | _033_;
  assign _039_ = _038_ ^ _037_;
  assign ctr_n[2] = down_i ? _039_ : _036_;
  assign _040_ = set_i ? val_i[3] : ctr_r[3];
  assign _041_ = _037_ & ~(_038_);
  assign _042_ = _041_ ^ _040_;
  assign ctr_n[3] = down_i ? _042_ : _040_;
  assign _043_ = set_i ? val_i[4] : ctr_r[4];
  assign _044_ = ~_043_;
  assign _045_ = _040_ | _036_;
  assign _046_ = _038_ & ~(_045_);
  assign _047_ = _046_ | _045_;
  assign _048_ = _047_ ^ _044_;
  assign ctr_n[4] = down_i ? _048_ : _043_;
  assign _049_ = set_i ? val_i[5] : ctr_r[5];
  assign _050_ = _044_ & ~(_047_);
  assign _051_ = _050_ ^ _049_;
  assign ctr_n[5] = down_i ? _051_ : _049_;
  assign _052_ = set_i ? val_i[6] : ctr_r[6];
  assign _053_ = ~_052_;
  assign _054_ = _049_ | _043_;
  assign _055_ = _047_ & ~(_054_);
  assign _056_ = _055_ | _054_;
  assign _057_ = _056_ ^ _053_;
  assign ctr_n[6] = down_i ? _057_ : _052_;
  assign _058_ = set_i ? val_i[7] : ctr_r[7];
  assign _059_ = _053_ & ~(_056_);
  assign _060_ = _059_ ^ _058_;
  assign ctr_n[7] = down_i ? _060_ : _058_;
  assign _061_ = set_i ? val_i[8] : ctr_r[8];
  assign _062_ = _058_ | _052_;
  assign _063_ = _054_ & ~(_062_);
  assign _064_ = _063_ | _062_;
  assign _065_ = _062_ | _054_;
  assign _066_ = _047_ & ~(_065_);
  assign _067_ = _066_ | _064_;
  assign _068_ = ~(_067_ ^ _061_);
  assign ctr_n[8] = down_i ? _068_ : _061_;
  assign _000_ = set_i ? val_i[9] : ctr_r[9];
  assign _001_ = ~(_067_ | _061_);
  assign _002_ = _001_ ^ _000_;
  assign ctr_n[9] = down_i ? _002_ : _000_;
  assign _003_ = set_i ? val_i[10] : ctr_r[10];
  assign _004_ = ~_003_;
  assign _005_ = _000_ | _061_;
  assign _006_ = _067_ & ~(_005_);
  assign _007_ = _006_ | _005_;
  assign _008_ = _007_ ^ _004_;
  assign ctr_n[10] = down_i ? _008_ : _003_;
  assign _009_ = set_i ? val_i[11] : ctr_r[11];
  assign _010_ = _004_ & ~(_007_);
  assign _011_ = _010_ ^ _009_;
  assign ctr_n[11] = down_i ? _011_ : _009_;
  assign _012_ = set_i ? val_i[12] : ctr_r[12];
  assign _013_ = _009_ | _003_;
  assign _014_ = _005_ & ~(_013_);
  assign _015_ = _014_ | _013_;
  assign _016_ = _013_ | _005_;
  assign _017_ = _067_ & ~(_016_);
  assign _018_ = _017_ | _015_;
  assign _019_ = ~(_018_ ^ _012_);
  assign ctr_n[12] = down_i ? _019_ : _012_;
  assign _020_ = set_i ? val_i[13] : ctr_r[13];
  assign _021_ = ~(_018_ | _012_);
  assign _022_ = _021_ ^ _020_;
  assign ctr_n[13] = down_i ? _022_ : _020_;
  assign _023_ = set_i ? val_i[14] : ctr_r[14];
  assign _024_ = ~_023_;
  assign _025_ = ~(_020_ | _012_);
  assign _026_ = _020_ | _012_;
  assign _027_ = _018_ & ~(_026_);
  assign _028_ = _027_ | ~(_025_);
  assign _029_ = _028_ ^ _024_;
  assign ctr_n[14] = down_i ? _029_ : _023_;
  assign _030_ = set_i ? val_i[15] : ctr_r[15];
  assign _031_ = _024_ & ~(_028_);
  assign _032_ = _031_ ^ _030_;
  assign ctr_n[15] = down_i ? _032_ : _030_;
  always @(posedge clk_i)
    if (reset_i) ctr_r[0] <= 1'h0;
    else ctr_r[0] <= ctr_n[0];
  always @(posedge clk_i)
    if (reset_i) ctr_r[1] <= 1'h0;
    else ctr_r[1] <= ctr_n[1];
  always @(posedge clk_i)
    if (reset_i) ctr_r[2] <= 1'h0;
    else ctr_r[2] <= ctr_n[2];
  always @(posedge clk_i)
    if (reset_i) ctr_r[3] <= 1'h0;
    else ctr_r[3] <= ctr_n[3];
  always @(posedge clk_i)
    if (reset_i) ctr_r[4] <= 1'h0;
    else ctr_r[4] <= ctr_n[4];
  always @(posedge clk_i)
    if (reset_i) ctr_r[5] <= 1'h0;
    else ctr_r[5] <= ctr_n[5];
  always @(posedge clk_i)
    if (reset_i) ctr_r[6] <= 1'h0;
    else ctr_r[6] <= ctr_n[6];
  always @(posedge clk_i)
    if (reset_i) ctr_r[7] <= 1'h0;
    else ctr_r[7] <= ctr_n[7];
  always @(posedge clk_i)
    if (reset_i) ctr_r[8] <= 1'h0;
    else ctr_r[8] <= ctr_n[8];
  always @(posedge clk_i)
    if (reset_i) ctr_r[9] <= 1'h0;
    else ctr_r[9] <= ctr_n[9];
  always @(posedge clk_i)
    if (reset_i) ctr_r[10] <= 1'h0;
    else ctr_r[10] <= ctr_n[10];
  always @(posedge clk_i)
    if (reset_i) ctr_r[11] <= 1'h0;
    else ctr_r[11] <= ctr_n[11];
  always @(posedge clk_i)
    if (reset_i) ctr_r[12] <= 1'h0;
    else ctr_r[12] <= ctr_n[12];
  always @(posedge clk_i)
    if (reset_i) ctr_r[13] <= 1'h0;
    else ctr_r[13] <= ctr_n[13];
  always @(posedge clk_i)
    if (reset_i) ctr_r[14] <= 1'h0;
    else ctr_r[14] <= ctr_n[14];
  always @(posedge clk_i)
    if (reset_i) ctr_r[15] <= 1'h0;
    else ctr_r[15] <= ctr_n[15];
  assign count_r_o = ctr_r;
endmodule
