module bsg_async_fifo(w_clk_i, w_reset_i, w_enq_i, w_data_i, w_full_o, r_clk_i, r_reset_i, r_deq_i, r_data_o, r_valid_o);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire [9:0] \MSYNC_1r1w.r_addr_i ;
  wire [15:0] \MSYNC_1r1w.r_data_o ;
  wire \MSYNC_1r1w.r_v_i ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[0] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1000] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1001] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1002] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1003] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1004] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1005] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1006] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1007] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1008] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1009] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[100] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1010] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1011] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1012] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1013] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1014] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1015] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1016] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1017] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1018] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1019] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[101] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1020] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1021] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1022] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1023] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[102] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[103] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[104] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[105] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[106] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[107] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[108] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[109] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[10] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[110] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[111] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[112] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[113] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[114] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[115] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[116] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[117] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[118] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[119] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[11] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[120] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[121] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[122] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[123] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[124] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[125] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[126] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[127] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[128] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[129] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[12] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[130] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[131] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[132] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[133] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[134] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[135] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[136] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[137] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[138] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[139] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[13] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[140] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[141] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[142] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[143] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[144] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[145] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[146] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[147] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[148] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[149] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[14] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[150] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[151] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[152] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[153] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[154] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[155] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[156] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[157] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[158] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[159] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[15] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[160] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[161] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[162] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[163] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[164] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[165] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[166] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[167] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[168] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[169] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[16] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[170] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[171] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[172] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[173] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[174] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[175] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[176] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[177] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[178] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[179] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[17] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[180] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[181] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[182] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[183] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[184] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[185] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[186] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[187] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[188] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[189] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[18] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[190] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[191] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[192] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[193] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[194] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[195] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[196] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[197] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[198] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[199] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[19] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[1] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[200] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[201] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[202] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[203] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[204] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[205] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[206] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[207] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[208] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[209] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[20] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[210] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[211] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[212] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[213] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[214] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[215] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[216] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[217] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[218] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[219] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[21] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[220] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[221] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[222] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[223] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[224] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[225] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[226] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[227] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[228] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[229] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[22] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[230] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[231] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[232] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[233] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[234] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[235] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[236] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[237] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[238] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[239] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[23] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[240] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[241] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[242] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[243] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[244] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[245] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[246] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[247] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[248] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[249] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[24] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[250] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[251] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[252] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[253] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[254] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[255] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[256] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[257] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[258] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[259] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[25] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[260] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[261] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[262] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[263] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[264] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[265] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[266] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[267] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[268] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[269] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[26] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[270] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[271] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[272] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[273] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[274] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[275] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[276] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[277] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[278] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[279] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[27] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[280] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[281] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[282] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[283] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[284] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[285] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[286] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[287] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[288] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[289] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[28] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[290] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[291] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[292] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[293] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[294] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[295] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[296] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[297] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[298] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[299] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[29] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[2] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[300] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[301] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[302] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[303] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[304] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[305] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[306] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[307] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[308] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[309] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[30] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[310] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[311] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[312] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[313] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[314] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[315] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[316] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[317] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[318] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[319] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[31] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[320] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[321] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[322] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[323] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[324] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[325] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[326] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[327] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[328] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[329] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[32] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[330] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[331] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[332] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[333] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[334] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[335] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[336] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[337] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[338] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[339] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[33] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[340] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[341] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[342] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[343] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[344] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[345] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[346] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[347] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[348] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[349] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[34] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[350] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[351] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[352] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[353] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[354] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[355] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[356] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[357] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[358] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[359] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[35] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[360] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[361] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[362] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[363] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[364] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[365] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[366] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[367] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[368] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[369] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[36] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[370] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[371] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[372] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[373] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[374] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[375] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[376] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[377] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[378] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[379] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[37] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[380] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[381] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[382] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[383] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[384] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[385] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[386] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[387] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[388] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[389] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[38] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[390] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[391] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[392] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[393] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[394] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[395] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[396] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[397] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[398] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[399] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[39] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[3] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[400] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[401] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[402] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[403] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[404] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[405] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[406] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[407] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[408] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[409] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[40] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[410] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[411] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[412] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[413] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[414] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[415] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[416] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[417] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[418] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[419] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[41] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[420] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[421] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[422] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[423] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[424] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[425] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[426] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[427] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[428] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[429] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[42] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[430] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[431] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[432] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[433] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[434] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[435] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[436] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[437] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[438] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[439] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[43] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[440] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[441] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[442] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[443] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[444] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[445] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[446] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[447] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[448] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[449] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[44] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[450] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[451] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[452] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[453] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[454] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[455] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[456] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[457] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[458] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[459] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[45] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[460] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[461] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[462] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[463] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[464] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[465] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[466] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[467] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[468] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[469] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[46] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[470] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[471] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[472] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[473] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[474] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[475] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[476] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[477] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[478] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[479] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[47] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[480] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[481] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[482] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[483] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[484] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[485] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[486] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[487] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[488] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[489] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[48] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[490] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[491] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[492] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[493] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[494] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[495] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[496] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[497] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[498] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[499] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[49] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[4] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[500] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[501] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[502] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[503] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[504] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[505] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[506] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[507] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[508] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[509] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[50] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[510] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[511] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[512] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[513] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[514] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[515] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[516] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[517] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[518] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[519] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[51] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[520] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[521] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[522] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[523] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[524] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[525] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[526] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[527] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[528] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[529] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[52] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[530] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[531] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[532] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[533] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[534] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[535] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[536] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[537] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[538] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[539] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[53] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[540] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[541] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[542] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[543] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[544] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[545] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[546] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[547] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[548] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[549] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[54] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[550] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[551] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[552] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[553] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[554] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[555] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[556] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[557] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[558] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[559] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[55] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[560] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[561] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[562] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[563] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[564] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[565] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[566] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[567] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[568] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[569] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[56] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[570] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[571] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[572] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[573] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[574] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[575] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[576] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[577] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[578] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[579] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[57] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[580] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[581] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[582] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[583] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[584] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[585] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[586] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[587] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[588] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[589] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[58] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[590] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[591] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[592] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[593] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[594] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[595] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[596] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[597] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[598] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[599] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[59] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[5] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[600] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[601] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[602] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[603] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[604] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[605] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[606] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[607] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[608] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[609] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[60] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[610] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[611] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[612] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[613] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[614] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[615] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[616] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[617] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[618] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[619] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[61] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[620] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[621] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[622] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[623] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[624] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[625] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[626] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[627] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[628] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[629] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[62] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[630] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[631] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[632] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[633] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[634] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[635] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[636] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[637] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[638] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[639] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[63] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[640] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[641] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[642] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[643] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[644] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[645] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[646] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[647] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[648] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[649] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[64] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[650] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[651] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[652] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[653] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[654] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[655] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[656] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[657] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[658] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[659] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[65] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[660] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[661] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[662] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[663] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[664] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[665] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[666] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[667] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[668] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[669] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[66] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[670] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[671] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[672] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[673] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[674] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[675] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[676] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[677] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[678] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[679] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[67] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[680] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[681] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[682] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[683] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[684] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[685] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[686] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[687] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[688] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[689] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[68] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[690] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[691] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[692] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[693] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[694] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[695] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[696] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[697] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[698] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[699] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[69] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[6] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[700] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[701] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[702] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[703] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[704] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[705] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[706] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[707] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[708] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[709] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[70] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[710] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[711] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[712] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[713] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[714] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[715] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[716] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[717] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[718] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[719] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[71] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[720] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[721] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[722] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[723] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[724] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[725] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[726] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[727] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[728] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[729] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[72] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[730] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[731] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[732] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[733] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[734] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[735] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[736] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[737] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[738] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[739] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[73] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[740] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[741] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[742] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[743] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[744] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[745] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[746] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[747] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[748] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[749] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[74] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[750] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[751] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[752] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[753] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[754] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[755] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[756] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[757] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[758] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[759] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[75] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[760] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[761] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[762] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[763] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[764] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[765] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[766] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[767] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[768] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[769] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[76] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[770] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[771] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[772] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[773] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[774] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[775] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[776] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[777] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[778] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[779] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[77] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[780] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[781] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[782] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[783] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[784] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[785] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[786] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[787] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[788] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[789] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[78] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[790] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[791] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[792] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[793] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[794] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[795] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[796] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[797] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[798] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[799] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[79] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[7] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[800] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[801] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[802] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[803] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[804] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[805] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[806] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[807] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[808] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[809] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[80] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[810] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[811] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[812] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[813] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[814] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[815] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[816] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[817] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[818] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[819] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[81] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[820] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[821] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[822] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[823] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[824] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[825] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[826] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[827] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[828] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[829] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[82] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[830] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[831] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[832] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[833] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[834] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[835] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[836] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[837] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[838] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[839] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[83] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[840] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[841] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[842] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[843] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[844] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[845] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[846] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[847] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[848] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[849] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[84] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[850] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[851] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[852] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[853] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[854] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[855] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[856] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[857] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[858] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[859] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[85] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[860] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[861] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[862] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[863] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[864] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[865] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[866] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[867] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[868] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[869] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[86] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[870] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[871] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[872] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[873] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[874] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[875] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[876] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[877] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[878] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[879] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[87] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[880] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[881] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[882] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[883] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[884] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[885] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[886] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[887] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[888] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[889] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[88] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[890] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[891] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[892] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[893] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[894] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[895] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[896] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[897] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[898] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[899] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[89] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[8] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[900] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[901] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[902] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[903] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[904] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[905] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[906] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[907] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[908] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[909] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[90] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[910] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[911] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[912] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[913] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[914] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[915] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[916] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[917] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[918] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[919] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[91] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[920] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[921] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[922] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[923] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[924] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[925] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[926] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[927] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[928] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[929] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[92] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[930] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[931] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[932] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[933] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[934] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[935] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[936] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[937] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[938] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[939] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[93] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[940] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[941] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[942] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[943] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[944] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[945] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[946] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[947] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[948] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[949] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[94] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[950] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[951] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[952] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[953] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[954] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[955] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[956] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[957] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[958] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[959] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[95] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[960] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[961] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[962] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[963] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[964] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[965] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[966] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[967] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[968] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[969] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[96] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[970] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[971] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[972] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[973] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[974] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[975] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[976] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[977] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[978] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[979] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[97] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[980] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[981] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[982] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[983] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[984] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[985] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[986] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[987] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[988] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[989] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[98] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[990] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[991] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[992] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[993] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[994] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[995] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[996] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[997] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[998] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[999] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[99] ;
  reg [15:0] \MSYNC_1r1w.synth.nz.mem[9] ;
  wire [9:0] \MSYNC_1r1w.synth.r_addr_i ;
  wire [15:0] \MSYNC_1r1w.synth.r_data_o ;
  wire \MSYNC_1r1w.synth.r_v_i ;
  wire \MSYNC_1r1w.synth.unused0 ;
  wire \MSYNC_1r1w.synth.unused1 ;
  wire [9:0] \MSYNC_1r1w.synth.w_addr_i ;
  wire \MSYNC_1r1w.synth.w_clk_i ;
  wire [15:0] \MSYNC_1r1w.synth.w_data_i ;
  wire \MSYNC_1r1w.synth.w_reset_i ;
  wire \MSYNC_1r1w.synth.w_v_i ;
  wire [9:0] \MSYNC_1r1w.w_addr_i ;
  wire \MSYNC_1r1w.w_clk_i ;
  wire [15:0] \MSYNC_1r1w.w_data_i ;
  wire \MSYNC_1r1w.w_reset_i ;
  wire \MSYNC_1r1w.w_v_i ;
  wire [10:0] \bapg_rd.ptr_sync.iclk_data_o ;
  wire \bapg_rd.ptr_sync.iclk_i ;
  wire \bapg_rd.ptr_sync.iclk_reset_i ;
  wire [10:0] \bapg_rd.ptr_sync.oclk_data_o ;
  wire \bapg_rd.ptr_sync.oclk_i ;
  reg [7:0] \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r ;
  reg [7:0] \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r ;
  wire [7:0] \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r ;
  wire [7:0] \bapg_rd.ptr_sync.sync.p.maxb[0].blss.iclk_data_o ;
  wire \bapg_rd.ptr_sync.sync.p.maxb[0].blss.iclk_i ;
  wire \bapg_rd.ptr_sync.sync.p.maxb[0].blss.iclk_reset_i ;
  wire [7:0] \bapg_rd.ptr_sync.sync.p.maxb[0].blss.oclk_data_o ;
  wire \bapg_rd.ptr_sync.sync.p.maxb[0].blss.oclk_i ;
  reg [2:0] \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r ;
  reg [2:0] \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  reg [2:0] \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  wire [2:0] \bapg_rd.ptr_sync.sync.p.z.blss.iclk_data_o ;
  wire \bapg_rd.ptr_sync.sync.p.z.blss.iclk_i ;
  wire \bapg_rd.ptr_sync.sync.p.z.blss.iclk_reset_i ;
  wire [2:0] \bapg_rd.ptr_sync.sync.p.z.blss.oclk_data_o ;
  wire \bapg_rd.ptr_sync.sync.p.z.blss.oclk_i ;
  wire \bapg_rd.r_clk_i ;
  wire \bapg_rd.w_clk_i ;
  wire \bapg_rd.w_inc_i ;
  wire [10:0] \bapg_rd.w_ptr_binary_r_o ;
  wire [10:0] \bapg_rd.w_ptr_gray_r ;
  wire [10:0] \bapg_rd.w_ptr_gray_r_o ;
  wire [10:0] \bapg_rd.w_ptr_gray_r_rsync ;
  wire [10:0] \bapg_rd.w_ptr_gray_r_rsync_o ;
  reg [10:0] \bapg_rd.w_ptr_p1_r ;
  wire [10:0] \bapg_rd.w_ptr_p2 ;
  wire [10:0] \bapg_rd.w_ptr_r ;
  wire \bapg_rd.w_reset_i ;
  wire [10:0] \bapg_wr.ptr_sync.iclk_data_o ;
  wire \bapg_wr.ptr_sync.iclk_i ;
  wire \bapg_wr.ptr_sync.iclk_reset_i ;
  wire [10:0] \bapg_wr.ptr_sync.oclk_data_o ;
  wire \bapg_wr.ptr_sync.oclk_i ;
  reg [7:0] \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r ;
  reg [7:0] \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r ;
  wire [7:0] \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r ;
  wire [7:0] \bapg_wr.ptr_sync.sync.p.maxb[0].blss.iclk_data_o ;
  wire \bapg_wr.ptr_sync.sync.p.maxb[0].blss.iclk_i ;
  wire \bapg_wr.ptr_sync.sync.p.maxb[0].blss.iclk_reset_i ;
  wire [7:0] \bapg_wr.ptr_sync.sync.p.maxb[0].blss.oclk_data_o ;
  wire \bapg_wr.ptr_sync.sync.p.maxb[0].blss.oclk_i ;
  reg [2:0] \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r ;
  reg [2:0] \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  reg [2:0] \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  wire [2:0] \bapg_wr.ptr_sync.sync.p.z.blss.iclk_data_o ;
  wire \bapg_wr.ptr_sync.sync.p.z.blss.iclk_i ;
  wire \bapg_wr.ptr_sync.sync.p.z.blss.iclk_reset_i ;
  wire [2:0] \bapg_wr.ptr_sync.sync.p.z.blss.oclk_data_o ;
  wire \bapg_wr.ptr_sync.sync.p.z.blss.oclk_i ;
  wire \bapg_wr.r_clk_i ;
  wire \bapg_wr.w_clk_i ;
  wire \bapg_wr.w_inc_i ;
  wire [10:0] \bapg_wr.w_ptr_binary_r_o ;
  wire [10:0] \bapg_wr.w_ptr_gray_r ;
  wire [10:0] \bapg_wr.w_ptr_gray_r_o ;
  wire [10:0] \bapg_wr.w_ptr_gray_r_rsync ;
  wire [10:0] \bapg_wr.w_ptr_gray_r_rsync_o ;
  reg [10:0] \bapg_wr.w_ptr_p1_r ;
  wire [10:0] \bapg_wr.w_ptr_p2 ;
  wire [10:0] \bapg_wr.w_ptr_r ;
  wire \bapg_wr.w_reset_i ;
  input r_clk_i;
  wire r_clk_i;
  output [15:0] r_data_o;
  wire [15:0] r_data_o;
  wire [15:0] r_data_o_tmp;
  input r_deq_i;
  wire r_deq_i;
  wire [10:0] r_ptr_binary_r;
  wire [10:0] r_ptr_gray_r;
  wire [10:0] r_ptr_gray_r_wsync;
  input r_reset_i;
  wire r_reset_i;
  output r_valid_o;
  wire r_valid_o;
  wire r_valid_o_tmp;
  input w_clk_i;
  wire w_clk_i;
  input [15:0] w_data_i;
  wire [15:0] w_data_i;
  input w_enq_i;
  wire w_enq_i;
  output w_full_o;
  wire w_full_o;
  wire [10:0] w_ptr_binary_r;
  wire [10:0] w_ptr_gray_r;
  wire [10:0] w_ptr_gray_r_rsync;
  input w_reset_i;
  wire w_reset_i;
  assign \bapg_wr.w_ptr_p2 [0] = ~\bapg_wr.w_ptr_p1_r [0];
  assign \bapg_rd.w_ptr_p2 [0] = ~\bapg_rd.w_ptr_p1_r [0];
  assign _01042_ = \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [0] ^ \bapg_rd.w_ptr_p1_r [1];
  assign _01043_ = \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [1] ^ \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [1];
  assign _01044_ = _01043_ | _01042_;
  assign _01045_ = \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [2] ^ \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [2];
  assign _01046_ = \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [3] ^ \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [3];
  assign _01047_ = _01046_ | _01045_;
  assign _01048_ = _01047_ | _01044_;
  assign _01049_ = \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [4] ^ \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [4];
  assign _01050_ = \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [5] ^ \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [5];
  assign _01051_ = _01050_ | _01049_;
  assign _01052_ = \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [6] ^ \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [6];
  assign _01053_ = \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [7] ^ \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7];
  assign _01054_ = _01053_ | _01052_;
  assign _01055_ = _01054_ | _01051_;
  assign _01056_ = _01055_ | _01048_;
  assign _01057_ = \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] ^ \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  assign _01058_ = \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] ^ \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1];
  assign _01059_ = _01058_ | _01057_;
  assign _01060_ = \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [2] ^ \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [2];
  assign _01061_ = _01060_ | _01059_;
  assign r_valid_o = _01061_ | _01056_;
  assign _01062_ = ~(\bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [0] ^ \bapg_wr.w_ptr_p1_r [1]);
  assign _01063_ = \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [1] ^ \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [1];
  assign _01064_ = _01062_ & ~(_01063_);
  assign _01065_ = \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [2] ^ \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [2];
  assign _01066_ = \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [3] ^ \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [3];
  assign _01067_ = _01066_ | _01065_;
  assign _01068_ = _01064_ & ~(_01067_);
  assign _01069_ = \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [4] ^ \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [4];
  assign _01070_ = \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [5] ^ \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [5];
  assign _01071_ = _01070_ | _01069_;
  assign _01072_ = \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [6] ^ \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [6];
  assign _01073_ = \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [7] ^ \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7];
  assign _01074_ = _01073_ | _01072_;
  assign _01075_ = _01074_ | _01071_;
  assign _01076_ = _01068_ & ~(_01075_);
  assign _01077_ = \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] ^ \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  assign _01078_ = ~(\bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] ^ \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1]);
  assign _01079_ = _01078_ | _01077_;
  assign _01080_ = ~(\bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [2] ^ \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [2]);
  assign _01081_ = _01080_ | _01079_;
  assign w_full_o = _01076_ & ~(_01081_);
  assign _01082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [0] : \MSYNC_1r1w.synth.nz.mem[0] [0];
  assign _01083_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [0] : \MSYNC_1r1w.synth.nz.mem[2] [0];
  assign _01084_ = \bapg_rd.w_ptr_r [1] ? _01083_ : _01082_;
  assign _01085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [0] : \MSYNC_1r1w.synth.nz.mem[4] [0];
  assign _01086_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [0] : \MSYNC_1r1w.synth.nz.mem[6] [0];
  assign _01087_ = \bapg_rd.w_ptr_r [1] ? _01086_ : _01085_;
  assign _01088_ = \bapg_rd.w_ptr_r [2] ? _01087_ : _01084_;
  assign _01089_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [0] : \MSYNC_1r1w.synth.nz.mem[8] [0];
  assign _01090_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [0] : \MSYNC_1r1w.synth.nz.mem[10] [0];
  assign _01091_ = \bapg_rd.w_ptr_r [1] ? _01090_ : _01089_;
  assign _01092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [0] : \MSYNC_1r1w.synth.nz.mem[12] [0];
  assign _01093_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [0] : \MSYNC_1r1w.synth.nz.mem[14] [0];
  assign _01094_ = \bapg_rd.w_ptr_r [1] ? _01093_ : _01092_;
  assign _01095_ = \bapg_rd.w_ptr_r [2] ? _01094_ : _01091_;
  assign _01096_ = \bapg_rd.w_ptr_r [3] ? _01095_ : _01088_;
  assign _01097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [0] : \MSYNC_1r1w.synth.nz.mem[16] [0];
  assign _01098_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [0] : \MSYNC_1r1w.synth.nz.mem[18] [0];
  assign _01099_ = \bapg_rd.w_ptr_r [1] ? _01098_ : _01097_;
  assign _01100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [0] : \MSYNC_1r1w.synth.nz.mem[20] [0];
  assign _01101_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [0] : \MSYNC_1r1w.synth.nz.mem[22] [0];
  assign _01102_ = \bapg_rd.w_ptr_r [1] ? _01101_ : _01100_;
  assign _01103_ = \bapg_rd.w_ptr_r [2] ? _01102_ : _01099_;
  assign _01104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [0] : \MSYNC_1r1w.synth.nz.mem[24] [0];
  assign _01105_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [0] : \MSYNC_1r1w.synth.nz.mem[26] [0];
  assign _01106_ = \bapg_rd.w_ptr_r [1] ? _01105_ : _01104_;
  assign _01107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [0] : \MSYNC_1r1w.synth.nz.mem[28] [0];
  assign _01108_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [0] : \MSYNC_1r1w.synth.nz.mem[30] [0];
  assign _01109_ = \bapg_rd.w_ptr_r [1] ? _01108_ : _01107_;
  assign _01110_ = \bapg_rd.w_ptr_r [2] ? _01109_ : _01106_;
  assign _01111_ = \bapg_rd.w_ptr_r [3] ? _01110_ : _01103_;
  assign _01112_ = \bapg_rd.w_ptr_r [4] ? _01111_ : _01096_;
  assign _01113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [0] : \MSYNC_1r1w.synth.nz.mem[32] [0];
  assign _01114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [0] : \MSYNC_1r1w.synth.nz.mem[34] [0];
  assign _01115_ = \bapg_rd.w_ptr_r [1] ? _01114_ : _01113_;
  assign _01116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [0] : \MSYNC_1r1w.synth.nz.mem[36] [0];
  assign _01117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [0] : \MSYNC_1r1w.synth.nz.mem[38] [0];
  assign _01118_ = \bapg_rd.w_ptr_r [1] ? _01117_ : _01116_;
  assign _01119_ = \bapg_rd.w_ptr_r [2] ? _01118_ : _01115_;
  assign _01120_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [0] : \MSYNC_1r1w.synth.nz.mem[40] [0];
  assign _01121_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [0] : \MSYNC_1r1w.synth.nz.mem[42] [0];
  assign _01122_ = \bapg_rd.w_ptr_r [1] ? _01121_ : _01120_;
  assign _01123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [0] : \MSYNC_1r1w.synth.nz.mem[44] [0];
  assign _01124_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [0] : \MSYNC_1r1w.synth.nz.mem[46] [0];
  assign _01125_ = \bapg_rd.w_ptr_r [1] ? _01124_ : _01123_;
  assign _01126_ = \bapg_rd.w_ptr_r [2] ? _01125_ : _01122_;
  assign _01127_ = \bapg_rd.w_ptr_r [3] ? _01126_ : _01119_;
  assign _01128_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [0] : \MSYNC_1r1w.synth.nz.mem[48] [0];
  assign _01129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [0] : \MSYNC_1r1w.synth.nz.mem[50] [0];
  assign _01130_ = \bapg_rd.w_ptr_r [1] ? _01129_ : _01128_;
  assign _01131_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [0] : \MSYNC_1r1w.synth.nz.mem[52] [0];
  assign _01132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [0] : \MSYNC_1r1w.synth.nz.mem[54] [0];
  assign _01133_ = \bapg_rd.w_ptr_r [1] ? _01132_ : _01131_;
  assign _01134_ = \bapg_rd.w_ptr_r [2] ? _01133_ : _01130_;
  assign _01135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [0] : \MSYNC_1r1w.synth.nz.mem[56] [0];
  assign _01136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [0] : \MSYNC_1r1w.synth.nz.mem[58] [0];
  assign _01137_ = \bapg_rd.w_ptr_r [1] ? _01136_ : _01135_;
  assign _01138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [0] : \MSYNC_1r1w.synth.nz.mem[60] [0];
  assign _01139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [0] : \MSYNC_1r1w.synth.nz.mem[62] [0];
  assign _01140_ = \bapg_rd.w_ptr_r [1] ? _01139_ : _01138_;
  assign _01141_ = \bapg_rd.w_ptr_r [2] ? _01140_ : _01137_;
  assign _01142_ = \bapg_rd.w_ptr_r [3] ? _01141_ : _01134_;
  assign _01143_ = \bapg_rd.w_ptr_r [4] ? _01142_ : _01127_;
  assign _01144_ = \bapg_rd.w_ptr_r [5] ? _01143_ : _01112_;
  assign _01145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [0] : \MSYNC_1r1w.synth.nz.mem[64] [0];
  assign _01146_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [0] : \MSYNC_1r1w.synth.nz.mem[66] [0];
  assign _01147_ = \bapg_rd.w_ptr_r [1] ? _01146_ : _01145_;
  assign _01148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [0] : \MSYNC_1r1w.synth.nz.mem[68] [0];
  assign _01149_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [0] : \MSYNC_1r1w.synth.nz.mem[70] [0];
  assign _01150_ = \bapg_rd.w_ptr_r [1] ? _01149_ : _01148_;
  assign _01151_ = \bapg_rd.w_ptr_r [2] ? _01150_ : _01147_;
  assign _01152_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [0] : \MSYNC_1r1w.synth.nz.mem[72] [0];
  assign _01153_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [0] : \MSYNC_1r1w.synth.nz.mem[74] [0];
  assign _01154_ = \bapg_rd.w_ptr_r [1] ? _01153_ : _01152_;
  assign _01155_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [0] : \MSYNC_1r1w.synth.nz.mem[76] [0];
  assign _01156_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [0] : \MSYNC_1r1w.synth.nz.mem[78] [0];
  assign _01157_ = \bapg_rd.w_ptr_r [1] ? _01156_ : _01155_;
  assign _01158_ = \bapg_rd.w_ptr_r [2] ? _01157_ : _01154_;
  assign _01159_ = \bapg_rd.w_ptr_r [3] ? _01158_ : _01151_;
  assign _01160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [0] : \MSYNC_1r1w.synth.nz.mem[80] [0];
  assign _01161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [0] : \MSYNC_1r1w.synth.nz.mem[82] [0];
  assign _01162_ = \bapg_rd.w_ptr_r [1] ? _01161_ : _01160_;
  assign _01163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [0] : \MSYNC_1r1w.synth.nz.mem[84] [0];
  assign _01164_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [0] : \MSYNC_1r1w.synth.nz.mem[86] [0];
  assign _01165_ = \bapg_rd.w_ptr_r [1] ? _01164_ : _01163_;
  assign _01166_ = \bapg_rd.w_ptr_r [2] ? _01165_ : _01162_;
  assign _01167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [0] : \MSYNC_1r1w.synth.nz.mem[88] [0];
  assign _01168_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [0] : \MSYNC_1r1w.synth.nz.mem[90] [0];
  assign _01169_ = \bapg_rd.w_ptr_r [1] ? _01168_ : _01167_;
  assign _01170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [0] : \MSYNC_1r1w.synth.nz.mem[92] [0];
  assign _01171_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [0] : \MSYNC_1r1w.synth.nz.mem[94] [0];
  assign _01172_ = \bapg_rd.w_ptr_r [1] ? _01171_ : _01170_;
  assign _01173_ = \bapg_rd.w_ptr_r [2] ? _01172_ : _01169_;
  assign _01174_ = \bapg_rd.w_ptr_r [3] ? _01173_ : _01166_;
  assign _01175_ = \bapg_rd.w_ptr_r [4] ? _01174_ : _01159_;
  assign _01176_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [0] : \MSYNC_1r1w.synth.nz.mem[96] [0];
  assign _01177_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [0] : \MSYNC_1r1w.synth.nz.mem[98] [0];
  assign _01178_ = \bapg_rd.w_ptr_r [1] ? _01177_ : _01176_;
  assign _01179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [0] : \MSYNC_1r1w.synth.nz.mem[100] [0];
  assign _01180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [0] : \MSYNC_1r1w.synth.nz.mem[102] [0];
  assign _01181_ = \bapg_rd.w_ptr_r [1] ? _01180_ : _01179_;
  assign _01182_ = \bapg_rd.w_ptr_r [2] ? _01181_ : _01178_;
  assign _01183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [0] : \MSYNC_1r1w.synth.nz.mem[104] [0];
  assign _01184_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [0] : \MSYNC_1r1w.synth.nz.mem[106] [0];
  assign _01185_ = \bapg_rd.w_ptr_r [1] ? _01184_ : _01183_;
  assign _01186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [0] : \MSYNC_1r1w.synth.nz.mem[108] [0];
  assign _01187_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [0] : \MSYNC_1r1w.synth.nz.mem[110] [0];
  assign _01188_ = \bapg_rd.w_ptr_r [1] ? _01187_ : _01186_;
  assign _01189_ = \bapg_rd.w_ptr_r [2] ? _01188_ : _01185_;
  assign _01190_ = \bapg_rd.w_ptr_r [3] ? _01189_ : _01182_;
  assign _01191_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [0] : \MSYNC_1r1w.synth.nz.mem[112] [0];
  assign _01192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [0] : \MSYNC_1r1w.synth.nz.mem[114] [0];
  assign _01193_ = \bapg_rd.w_ptr_r [1] ? _01192_ : _01191_;
  assign _01194_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [0] : \MSYNC_1r1w.synth.nz.mem[116] [0];
  assign _01195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [0] : \MSYNC_1r1w.synth.nz.mem[118] [0];
  assign _01196_ = \bapg_rd.w_ptr_r [1] ? _01195_ : _01194_;
  assign _01197_ = \bapg_rd.w_ptr_r [2] ? _01196_ : _01193_;
  assign _01198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [0] : \MSYNC_1r1w.synth.nz.mem[120] [0];
  assign _01199_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [0] : \MSYNC_1r1w.synth.nz.mem[122] [0];
  assign _01200_ = \bapg_rd.w_ptr_r [1] ? _01199_ : _01198_;
  assign _01201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [0] : \MSYNC_1r1w.synth.nz.mem[124] [0];
  assign _01202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [0] : \MSYNC_1r1w.synth.nz.mem[126] [0];
  assign _01203_ = \bapg_rd.w_ptr_r [1] ? _01202_ : _01201_;
  assign _01204_ = \bapg_rd.w_ptr_r [2] ? _01203_ : _01200_;
  assign _01205_ = \bapg_rd.w_ptr_r [3] ? _01204_ : _01197_;
  assign _01206_ = \bapg_rd.w_ptr_r [4] ? _01205_ : _01190_;
  assign _01207_ = \bapg_rd.w_ptr_r [5] ? _01206_ : _01175_;
  assign _01208_ = \bapg_rd.w_ptr_r [6] ? _01207_ : _01144_;
  assign _01209_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [0] : \MSYNC_1r1w.synth.nz.mem[128] [0];
  assign _01210_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [0] : \MSYNC_1r1w.synth.nz.mem[130] [0];
  assign _01211_ = \bapg_rd.w_ptr_r [1] ? _01210_ : _01209_;
  assign _01212_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [0] : \MSYNC_1r1w.synth.nz.mem[132] [0];
  assign _01213_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [0] : \MSYNC_1r1w.synth.nz.mem[134] [0];
  assign _01214_ = \bapg_rd.w_ptr_r [1] ? _01213_ : _01212_;
  assign _01215_ = \bapg_rd.w_ptr_r [2] ? _01214_ : _01211_;
  assign _01216_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [0] : \MSYNC_1r1w.synth.nz.mem[136] [0];
  assign _01217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [0] : \MSYNC_1r1w.synth.nz.mem[138] [0];
  assign _01218_ = \bapg_rd.w_ptr_r [1] ? _01217_ : _01216_;
  assign _01219_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [0] : \MSYNC_1r1w.synth.nz.mem[140] [0];
  assign _01220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [0] : \MSYNC_1r1w.synth.nz.mem[142] [0];
  assign _01221_ = \bapg_rd.w_ptr_r [1] ? _01220_ : _01219_;
  assign _01222_ = \bapg_rd.w_ptr_r [2] ? _01221_ : _01218_;
  assign _01223_ = \bapg_rd.w_ptr_r [3] ? _01222_ : _01215_;
  assign _01224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [0] : \MSYNC_1r1w.synth.nz.mem[144] [0];
  assign _01225_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [0] : \MSYNC_1r1w.synth.nz.mem[146] [0];
  assign _01226_ = \bapg_rd.w_ptr_r [1] ? _01225_ : _01224_;
  assign _01227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [0] : \MSYNC_1r1w.synth.nz.mem[148] [0];
  assign _01228_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [0] : \MSYNC_1r1w.synth.nz.mem[150] [0];
  assign _01229_ = \bapg_rd.w_ptr_r [1] ? _01228_ : _01227_;
  assign _01230_ = \bapg_rd.w_ptr_r [2] ? _01229_ : _01226_;
  assign _01231_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [0] : \MSYNC_1r1w.synth.nz.mem[152] [0];
  assign _01232_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [0] : \MSYNC_1r1w.synth.nz.mem[154] [0];
  assign _01233_ = \bapg_rd.w_ptr_r [1] ? _01232_ : _01231_;
  assign _01234_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [0] : \MSYNC_1r1w.synth.nz.mem[156] [0];
  assign _01235_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [0] : \MSYNC_1r1w.synth.nz.mem[158] [0];
  assign _01236_ = \bapg_rd.w_ptr_r [1] ? _01235_ : _01234_;
  assign _01237_ = \bapg_rd.w_ptr_r [2] ? _01236_ : _01233_;
  assign _01238_ = \bapg_rd.w_ptr_r [3] ? _01237_ : _01230_;
  assign _01239_ = \bapg_rd.w_ptr_r [4] ? _01238_ : _01223_;
  assign _01240_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [0] : \MSYNC_1r1w.synth.nz.mem[160] [0];
  assign _01241_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [0] : \MSYNC_1r1w.synth.nz.mem[162] [0];
  assign _01242_ = \bapg_rd.w_ptr_r [1] ? _01241_ : _01240_;
  assign _01243_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [0] : \MSYNC_1r1w.synth.nz.mem[164] [0];
  assign _01244_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [0] : \MSYNC_1r1w.synth.nz.mem[166] [0];
  assign _01245_ = \bapg_rd.w_ptr_r [1] ? _01244_ : _01243_;
  assign _01246_ = \bapg_rd.w_ptr_r [2] ? _01245_ : _01242_;
  assign _01247_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [0] : \MSYNC_1r1w.synth.nz.mem[168] [0];
  assign _01248_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [0] : \MSYNC_1r1w.synth.nz.mem[170] [0];
  assign _01249_ = \bapg_rd.w_ptr_r [1] ? _01248_ : _01247_;
  assign _01250_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [0] : \MSYNC_1r1w.synth.nz.mem[172] [0];
  assign _01251_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [0] : \MSYNC_1r1w.synth.nz.mem[174] [0];
  assign _01252_ = \bapg_rd.w_ptr_r [1] ? _01251_ : _01250_;
  assign _01253_ = \bapg_rd.w_ptr_r [2] ? _01252_ : _01249_;
  assign _01254_ = \bapg_rd.w_ptr_r [3] ? _01253_ : _01246_;
  assign _01255_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [0] : \MSYNC_1r1w.synth.nz.mem[176] [0];
  assign _01256_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [0] : \MSYNC_1r1w.synth.nz.mem[178] [0];
  assign _01257_ = \bapg_rd.w_ptr_r [1] ? _01256_ : _01255_;
  assign _01258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [0] : \MSYNC_1r1w.synth.nz.mem[180] [0];
  assign _01259_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [0] : \MSYNC_1r1w.synth.nz.mem[182] [0];
  assign _01260_ = \bapg_rd.w_ptr_r [1] ? _01259_ : _01258_;
  assign _01261_ = \bapg_rd.w_ptr_r [2] ? _01260_ : _01257_;
  assign _01262_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [0] : \MSYNC_1r1w.synth.nz.mem[184] [0];
  assign _01263_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [0] : \MSYNC_1r1w.synth.nz.mem[186] [0];
  assign _01264_ = \bapg_rd.w_ptr_r [1] ? _01263_ : _01262_;
  assign _01265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [0] : \MSYNC_1r1w.synth.nz.mem[188] [0];
  assign _01266_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [0] : \MSYNC_1r1w.synth.nz.mem[190] [0];
  assign _01267_ = \bapg_rd.w_ptr_r [1] ? _01266_ : _01265_;
  assign _01268_ = \bapg_rd.w_ptr_r [2] ? _01267_ : _01264_;
  assign _01269_ = \bapg_rd.w_ptr_r [3] ? _01268_ : _01261_;
  assign _01270_ = \bapg_rd.w_ptr_r [4] ? _01269_ : _01254_;
  assign _01271_ = \bapg_rd.w_ptr_r [5] ? _01270_ : _01239_;
  assign _01272_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [0] : \MSYNC_1r1w.synth.nz.mem[192] [0];
  assign _01273_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [0] : \MSYNC_1r1w.synth.nz.mem[194] [0];
  assign _01274_ = \bapg_rd.w_ptr_r [1] ? _01273_ : _01272_;
  assign _01275_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [0] : \MSYNC_1r1w.synth.nz.mem[196] [0];
  assign _01276_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [0] : \MSYNC_1r1w.synth.nz.mem[198] [0];
  assign _01277_ = \bapg_rd.w_ptr_r [1] ? _01276_ : _01275_;
  assign _01278_ = \bapg_rd.w_ptr_r [2] ? _01277_ : _01274_;
  assign _01279_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [0] : \MSYNC_1r1w.synth.nz.mem[200] [0];
  assign _01280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [0] : \MSYNC_1r1w.synth.nz.mem[202] [0];
  assign _01281_ = \bapg_rd.w_ptr_r [1] ? _01280_ : _01279_;
  assign _01282_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [0] : \MSYNC_1r1w.synth.nz.mem[204] [0];
  assign _01283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [0] : \MSYNC_1r1w.synth.nz.mem[206] [0];
  assign _01284_ = \bapg_rd.w_ptr_r [1] ? _01283_ : _01282_;
  assign _01285_ = \bapg_rd.w_ptr_r [2] ? _01284_ : _01281_;
  assign _01286_ = \bapg_rd.w_ptr_r [3] ? _01285_ : _01278_;
  assign _01287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [0] : \MSYNC_1r1w.synth.nz.mem[208] [0];
  assign _01288_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [0] : \MSYNC_1r1w.synth.nz.mem[210] [0];
  assign _01289_ = \bapg_rd.w_ptr_r [1] ? _01288_ : _01287_;
  assign _01290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [0] : \MSYNC_1r1w.synth.nz.mem[212] [0];
  assign _01291_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [0] : \MSYNC_1r1w.synth.nz.mem[214] [0];
  assign _01292_ = \bapg_rd.w_ptr_r [1] ? _01291_ : _01290_;
  assign _01293_ = \bapg_rd.w_ptr_r [2] ? _01292_ : _01289_;
  assign _01294_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [0] : \MSYNC_1r1w.synth.nz.mem[216] [0];
  assign _01295_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [0] : \MSYNC_1r1w.synth.nz.mem[218] [0];
  assign _01296_ = \bapg_rd.w_ptr_r [1] ? _01295_ : _01294_;
  assign _01297_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [0] : \MSYNC_1r1w.synth.nz.mem[220] [0];
  assign _01298_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [0] : \MSYNC_1r1w.synth.nz.mem[222] [0];
  assign _01299_ = \bapg_rd.w_ptr_r [1] ? _01298_ : _01297_;
  assign _01300_ = \bapg_rd.w_ptr_r [2] ? _01299_ : _01296_;
  assign _01301_ = \bapg_rd.w_ptr_r [3] ? _01300_ : _01293_;
  assign _01302_ = \bapg_rd.w_ptr_r [4] ? _01301_ : _01286_;
  assign _01303_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [0] : \MSYNC_1r1w.synth.nz.mem[224] [0];
  assign _01304_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [0] : \MSYNC_1r1w.synth.nz.mem[226] [0];
  assign _01305_ = \bapg_rd.w_ptr_r [1] ? _01304_ : _01303_;
  assign _01306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [0] : \MSYNC_1r1w.synth.nz.mem[228] [0];
  assign _01307_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [0] : \MSYNC_1r1w.synth.nz.mem[230] [0];
  assign _01308_ = \bapg_rd.w_ptr_r [1] ? _01307_ : _01306_;
  assign _01309_ = \bapg_rd.w_ptr_r [2] ? _01308_ : _01305_;
  assign _01310_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [0] : \MSYNC_1r1w.synth.nz.mem[232] [0];
  assign _01311_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [0] : \MSYNC_1r1w.synth.nz.mem[234] [0];
  assign _01312_ = \bapg_rd.w_ptr_r [1] ? _01311_ : _01310_;
  assign _01313_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [0] : \MSYNC_1r1w.synth.nz.mem[236] [0];
  assign _01314_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [0] : \MSYNC_1r1w.synth.nz.mem[238] [0];
  assign _01315_ = \bapg_rd.w_ptr_r [1] ? _01314_ : _01313_;
  assign _01316_ = \bapg_rd.w_ptr_r [2] ? _01315_ : _01312_;
  assign _01317_ = \bapg_rd.w_ptr_r [3] ? _01316_ : _01309_;
  assign _01318_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [0] : \MSYNC_1r1w.synth.nz.mem[240] [0];
  assign _01319_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [0] : \MSYNC_1r1w.synth.nz.mem[242] [0];
  assign _01320_ = \bapg_rd.w_ptr_r [1] ? _01319_ : _01318_;
  assign _01321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [0] : \MSYNC_1r1w.synth.nz.mem[244] [0];
  assign _01322_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [0] : \MSYNC_1r1w.synth.nz.mem[246] [0];
  assign _01323_ = \bapg_rd.w_ptr_r [1] ? _01322_ : _01321_;
  assign _01324_ = \bapg_rd.w_ptr_r [2] ? _01323_ : _01320_;
  assign _01325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [0] : \MSYNC_1r1w.synth.nz.mem[248] [0];
  assign _01326_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [0] : \MSYNC_1r1w.synth.nz.mem[250] [0];
  assign _01327_ = \bapg_rd.w_ptr_r [1] ? _01326_ : _01325_;
  assign _01328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [0] : \MSYNC_1r1w.synth.nz.mem[252] [0];
  assign _01329_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [0] : \MSYNC_1r1w.synth.nz.mem[254] [0];
  assign _01330_ = \bapg_rd.w_ptr_r [1] ? _01329_ : _01328_;
  assign _01331_ = \bapg_rd.w_ptr_r [2] ? _01330_ : _01327_;
  assign _01332_ = \bapg_rd.w_ptr_r [3] ? _01331_ : _01324_;
  assign _01333_ = \bapg_rd.w_ptr_r [4] ? _01332_ : _01317_;
  assign _01334_ = \bapg_rd.w_ptr_r [5] ? _01333_ : _01302_;
  assign _01335_ = \bapg_rd.w_ptr_r [6] ? _01334_ : _01271_;
  assign _01336_ = \bapg_rd.w_ptr_r [7] ? _01335_ : _01208_;
  assign _01337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [0] : \MSYNC_1r1w.synth.nz.mem[256] [0];
  assign _01338_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [0] : \MSYNC_1r1w.synth.nz.mem[258] [0];
  assign _01339_ = \bapg_rd.w_ptr_r [1] ? _01338_ : _01337_;
  assign _01340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [0] : \MSYNC_1r1w.synth.nz.mem[260] [0];
  assign _01341_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [0] : \MSYNC_1r1w.synth.nz.mem[262] [0];
  assign _01342_ = \bapg_rd.w_ptr_r [1] ? _01341_ : _01340_;
  assign _01343_ = \bapg_rd.w_ptr_r [2] ? _01342_ : _01339_;
  assign _01344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [0] : \MSYNC_1r1w.synth.nz.mem[264] [0];
  assign _01345_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [0] : \MSYNC_1r1w.synth.nz.mem[266] [0];
  assign _01346_ = \bapg_rd.w_ptr_r [1] ? _01345_ : _01344_;
  assign _01347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [0] : \MSYNC_1r1w.synth.nz.mem[268] [0];
  assign _01348_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [0] : \MSYNC_1r1w.synth.nz.mem[270] [0];
  assign _01349_ = \bapg_rd.w_ptr_r [1] ? _01348_ : _01347_;
  assign _01350_ = \bapg_rd.w_ptr_r [2] ? _01349_ : _01346_;
  assign _01351_ = \bapg_rd.w_ptr_r [3] ? _01350_ : _01343_;
  assign _01352_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [0] : \MSYNC_1r1w.synth.nz.mem[272] [0];
  assign _01353_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [0] : \MSYNC_1r1w.synth.nz.mem[274] [0];
  assign _01354_ = \bapg_rd.w_ptr_r [1] ? _01353_ : _01352_;
  assign _01355_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [0] : \MSYNC_1r1w.synth.nz.mem[276] [0];
  assign _01356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [0] : \MSYNC_1r1w.synth.nz.mem[278] [0];
  assign _01357_ = \bapg_rd.w_ptr_r [1] ? _01356_ : _01355_;
  assign _01358_ = \bapg_rd.w_ptr_r [2] ? _01357_ : _01354_;
  assign _01359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [0] : \MSYNC_1r1w.synth.nz.mem[280] [0];
  assign _01360_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [0] : \MSYNC_1r1w.synth.nz.mem[282] [0];
  assign _01361_ = \bapg_rd.w_ptr_r [1] ? _01360_ : _01359_;
  assign _01362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [0] : \MSYNC_1r1w.synth.nz.mem[284] [0];
  assign _01363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [0] : \MSYNC_1r1w.synth.nz.mem[286] [0];
  assign _01364_ = \bapg_rd.w_ptr_r [1] ? _01363_ : _01362_;
  assign _01365_ = \bapg_rd.w_ptr_r [2] ? _01364_ : _01361_;
  assign _01366_ = \bapg_rd.w_ptr_r [3] ? _01365_ : _01358_;
  assign _01367_ = \bapg_rd.w_ptr_r [4] ? _01366_ : _01351_;
  assign _01368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [0] : \MSYNC_1r1w.synth.nz.mem[288] [0];
  assign _01369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [0] : \MSYNC_1r1w.synth.nz.mem[290] [0];
  assign _01370_ = \bapg_rd.w_ptr_r [1] ? _01369_ : _01368_;
  assign _01371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [0] : \MSYNC_1r1w.synth.nz.mem[292] [0];
  assign _01372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [0] : \MSYNC_1r1w.synth.nz.mem[294] [0];
  assign _01373_ = \bapg_rd.w_ptr_r [1] ? _01372_ : _01371_;
  assign _01374_ = \bapg_rd.w_ptr_r [2] ? _01373_ : _01370_;
  assign _01375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [0] : \MSYNC_1r1w.synth.nz.mem[296] [0];
  assign _01376_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [0] : \MSYNC_1r1w.synth.nz.mem[298] [0];
  assign _01377_ = \bapg_rd.w_ptr_r [1] ? _01376_ : _01375_;
  assign _01378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [0] : \MSYNC_1r1w.synth.nz.mem[300] [0];
  assign _01379_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [0] : \MSYNC_1r1w.synth.nz.mem[302] [0];
  assign _01380_ = \bapg_rd.w_ptr_r [1] ? _01379_ : _01378_;
  assign _01381_ = \bapg_rd.w_ptr_r [2] ? _01380_ : _01377_;
  assign _01382_ = \bapg_rd.w_ptr_r [3] ? _01381_ : _01374_;
  assign _01383_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [0] : \MSYNC_1r1w.synth.nz.mem[304] [0];
  assign _01384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [0] : \MSYNC_1r1w.synth.nz.mem[306] [0];
  assign _01385_ = \bapg_rd.w_ptr_r [1] ? _01384_ : _01383_;
  assign _01386_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [0] : \MSYNC_1r1w.synth.nz.mem[308] [0];
  assign _01387_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [0] : \MSYNC_1r1w.synth.nz.mem[310] [0];
  assign _01388_ = \bapg_rd.w_ptr_r [1] ? _01387_ : _01386_;
  assign _01389_ = \bapg_rd.w_ptr_r [2] ? _01388_ : _01385_;
  assign _01390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [0] : \MSYNC_1r1w.synth.nz.mem[312] [0];
  assign _01391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [0] : \MSYNC_1r1w.synth.nz.mem[314] [0];
  assign _01392_ = \bapg_rd.w_ptr_r [1] ? _01391_ : _01390_;
  assign _01393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [0] : \MSYNC_1r1w.synth.nz.mem[316] [0];
  assign _01394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [0] : \MSYNC_1r1w.synth.nz.mem[318] [0];
  assign _01395_ = \bapg_rd.w_ptr_r [1] ? _01394_ : _01393_;
  assign _01396_ = \bapg_rd.w_ptr_r [2] ? _01395_ : _01392_;
  assign _01397_ = \bapg_rd.w_ptr_r [3] ? _01396_ : _01389_;
  assign _01398_ = \bapg_rd.w_ptr_r [4] ? _01397_ : _01382_;
  assign _01399_ = \bapg_rd.w_ptr_r [5] ? _01398_ : _01367_;
  assign _01400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [0] : \MSYNC_1r1w.synth.nz.mem[320] [0];
  assign _01401_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [0] : \MSYNC_1r1w.synth.nz.mem[322] [0];
  assign _01402_ = \bapg_rd.w_ptr_r [1] ? _01401_ : _01400_;
  assign _01403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [0] : \MSYNC_1r1w.synth.nz.mem[324] [0];
  assign _01404_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [0] : \MSYNC_1r1w.synth.nz.mem[326] [0];
  assign _01405_ = \bapg_rd.w_ptr_r [1] ? _01404_ : _01403_;
  assign _01406_ = \bapg_rd.w_ptr_r [2] ? _01405_ : _01402_;
  assign _01407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [0] : \MSYNC_1r1w.synth.nz.mem[328] [0];
  assign _01408_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [0] : \MSYNC_1r1w.synth.nz.mem[330] [0];
  assign _01409_ = \bapg_rd.w_ptr_r [1] ? _01408_ : _01407_;
  assign _01410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [0] : \MSYNC_1r1w.synth.nz.mem[332] [0];
  assign _01411_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [0] : \MSYNC_1r1w.synth.nz.mem[334] [0];
  assign _01412_ = \bapg_rd.w_ptr_r [1] ? _01411_ : _01410_;
  assign _01413_ = \bapg_rd.w_ptr_r [2] ? _01412_ : _01409_;
  assign _01414_ = \bapg_rd.w_ptr_r [3] ? _01413_ : _01406_;
  assign _01415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [0] : \MSYNC_1r1w.synth.nz.mem[336] [0];
  assign _01416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [0] : \MSYNC_1r1w.synth.nz.mem[338] [0];
  assign _01417_ = \bapg_rd.w_ptr_r [1] ? _01416_ : _01415_;
  assign _01418_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [0] : \MSYNC_1r1w.synth.nz.mem[340] [0];
  assign _01419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [0] : \MSYNC_1r1w.synth.nz.mem[342] [0];
  assign _01420_ = \bapg_rd.w_ptr_r [1] ? _01419_ : _01418_;
  assign _01421_ = \bapg_rd.w_ptr_r [2] ? _01420_ : _01417_;
  assign _01422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [0] : \MSYNC_1r1w.synth.nz.mem[344] [0];
  assign _01423_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [0] : \MSYNC_1r1w.synth.nz.mem[346] [0];
  assign _01424_ = \bapg_rd.w_ptr_r [1] ? _01423_ : _01422_;
  assign _01425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [0] : \MSYNC_1r1w.synth.nz.mem[348] [0];
  assign _01426_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [0] : \MSYNC_1r1w.synth.nz.mem[350] [0];
  assign _01427_ = \bapg_rd.w_ptr_r [1] ? _01426_ : _01425_;
  assign _01428_ = \bapg_rd.w_ptr_r [2] ? _01427_ : _01424_;
  assign _01429_ = \bapg_rd.w_ptr_r [3] ? _01428_ : _01421_;
  assign _01430_ = \bapg_rd.w_ptr_r [4] ? _01429_ : _01414_;
  assign _01431_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [0] : \MSYNC_1r1w.synth.nz.mem[352] [0];
  assign _01432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [0] : \MSYNC_1r1w.synth.nz.mem[354] [0];
  assign _01433_ = \bapg_rd.w_ptr_r [1] ? _01432_ : _01431_;
  assign _01434_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [0] : \MSYNC_1r1w.synth.nz.mem[356] [0];
  assign _01435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [0] : \MSYNC_1r1w.synth.nz.mem[358] [0];
  assign _01436_ = \bapg_rd.w_ptr_r [1] ? _01435_ : _01434_;
  assign _01437_ = \bapg_rd.w_ptr_r [2] ? _01436_ : _01433_;
  assign _01438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [0] : \MSYNC_1r1w.synth.nz.mem[360] [0];
  assign _01439_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [0] : \MSYNC_1r1w.synth.nz.mem[362] [0];
  assign _01440_ = \bapg_rd.w_ptr_r [1] ? _01439_ : _01438_;
  assign _01441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [0] : \MSYNC_1r1w.synth.nz.mem[364] [0];
  assign _01442_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [0] : \MSYNC_1r1w.synth.nz.mem[366] [0];
  assign _01443_ = \bapg_rd.w_ptr_r [1] ? _01442_ : _01441_;
  assign _01444_ = \bapg_rd.w_ptr_r [2] ? _01443_ : _01440_;
  assign _01445_ = \bapg_rd.w_ptr_r [3] ? _01444_ : _01437_;
  assign _01446_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [0] : \MSYNC_1r1w.synth.nz.mem[368] [0];
  assign _01447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [0] : \MSYNC_1r1w.synth.nz.mem[370] [0];
  assign _01448_ = \bapg_rd.w_ptr_r [1] ? _01447_ : _01446_;
  assign _01449_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [0] : \MSYNC_1r1w.synth.nz.mem[372] [0];
  assign _01450_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [0] : \MSYNC_1r1w.synth.nz.mem[374] [0];
  assign _01451_ = \bapg_rd.w_ptr_r [1] ? _01450_ : _01449_;
  assign _01452_ = \bapg_rd.w_ptr_r [2] ? _01451_ : _01448_;
  assign _01453_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [0] : \MSYNC_1r1w.synth.nz.mem[376] [0];
  assign _01454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [0] : \MSYNC_1r1w.synth.nz.mem[378] [0];
  assign _01455_ = \bapg_rd.w_ptr_r [1] ? _01454_ : _01453_;
  assign _01456_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [0] : \MSYNC_1r1w.synth.nz.mem[380] [0];
  assign _01457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [0] : \MSYNC_1r1w.synth.nz.mem[382] [0];
  assign _01458_ = \bapg_rd.w_ptr_r [1] ? _01457_ : _01456_;
  assign _01459_ = \bapg_rd.w_ptr_r [2] ? _01458_ : _01455_;
  assign _01460_ = \bapg_rd.w_ptr_r [3] ? _01459_ : _01452_;
  assign _01461_ = \bapg_rd.w_ptr_r [4] ? _01460_ : _01445_;
  assign _01462_ = \bapg_rd.w_ptr_r [5] ? _01461_ : _01430_;
  assign _01463_ = \bapg_rd.w_ptr_r [6] ? _01462_ : _01399_;
  assign _01464_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [0] : \MSYNC_1r1w.synth.nz.mem[384] [0];
  assign _01465_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [0] : \MSYNC_1r1w.synth.nz.mem[386] [0];
  assign _01466_ = \bapg_rd.w_ptr_r [1] ? _01465_ : _01464_;
  assign _01467_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [0] : \MSYNC_1r1w.synth.nz.mem[388] [0];
  assign _01468_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [0] : \MSYNC_1r1w.synth.nz.mem[390] [0];
  assign _01469_ = \bapg_rd.w_ptr_r [1] ? _01468_ : _01467_;
  assign _01470_ = \bapg_rd.w_ptr_r [2] ? _01469_ : _01466_;
  assign _01471_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [0] : \MSYNC_1r1w.synth.nz.mem[392] [0];
  assign _01472_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [0] : \MSYNC_1r1w.synth.nz.mem[394] [0];
  assign _01473_ = \bapg_rd.w_ptr_r [1] ? _01472_ : _01471_;
  assign _01474_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [0] : \MSYNC_1r1w.synth.nz.mem[396] [0];
  assign _01475_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [0] : \MSYNC_1r1w.synth.nz.mem[398] [0];
  assign _01476_ = \bapg_rd.w_ptr_r [1] ? _01475_ : _01474_;
  assign _01477_ = \bapg_rd.w_ptr_r [2] ? _01476_ : _01473_;
  assign _01478_ = \bapg_rd.w_ptr_r [3] ? _01477_ : _01470_;
  assign _01479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [0] : \MSYNC_1r1w.synth.nz.mem[400] [0];
  assign _01480_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [0] : \MSYNC_1r1w.synth.nz.mem[402] [0];
  assign _01481_ = \bapg_rd.w_ptr_r [1] ? _01480_ : _01479_;
  assign _01482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [0] : \MSYNC_1r1w.synth.nz.mem[404] [0];
  assign _01483_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [0] : \MSYNC_1r1w.synth.nz.mem[406] [0];
  assign _01484_ = \bapg_rd.w_ptr_r [1] ? _01483_ : _01482_;
  assign _01485_ = \bapg_rd.w_ptr_r [2] ? _01484_ : _01481_;
  assign _01486_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [0] : \MSYNC_1r1w.synth.nz.mem[408] [0];
  assign _01487_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [0] : \MSYNC_1r1w.synth.nz.mem[410] [0];
  assign _01488_ = \bapg_rd.w_ptr_r [1] ? _01487_ : _01486_;
  assign _01489_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [0] : \MSYNC_1r1w.synth.nz.mem[412] [0];
  assign _01490_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [0] : \MSYNC_1r1w.synth.nz.mem[414] [0];
  assign _01491_ = \bapg_rd.w_ptr_r [1] ? _01490_ : _01489_;
  assign _01492_ = \bapg_rd.w_ptr_r [2] ? _01491_ : _01488_;
  assign _01493_ = \bapg_rd.w_ptr_r [3] ? _01492_ : _01485_;
  assign _01494_ = \bapg_rd.w_ptr_r [4] ? _01493_ : _01478_;
  assign _01495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [0] : \MSYNC_1r1w.synth.nz.mem[416] [0];
  assign _01496_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [0] : \MSYNC_1r1w.synth.nz.mem[418] [0];
  assign _01497_ = \bapg_rd.w_ptr_r [1] ? _01496_ : _01495_;
  assign _01498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [0] : \MSYNC_1r1w.synth.nz.mem[420] [0];
  assign _01499_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [0] : \MSYNC_1r1w.synth.nz.mem[422] [0];
  assign _01500_ = \bapg_rd.w_ptr_r [1] ? _01499_ : _01498_;
  assign _01501_ = \bapg_rd.w_ptr_r [2] ? _01500_ : _01497_;
  assign _01502_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [0] : \MSYNC_1r1w.synth.nz.mem[424] [0];
  assign _01503_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [0] : \MSYNC_1r1w.synth.nz.mem[426] [0];
  assign _01504_ = \bapg_rd.w_ptr_r [1] ? _01503_ : _01502_;
  assign _01505_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [0] : \MSYNC_1r1w.synth.nz.mem[428] [0];
  assign _01506_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [0] : \MSYNC_1r1w.synth.nz.mem[430] [0];
  assign _01507_ = \bapg_rd.w_ptr_r [1] ? _01506_ : _01505_;
  assign _01508_ = \bapg_rd.w_ptr_r [2] ? _01507_ : _01504_;
  assign _01509_ = \bapg_rd.w_ptr_r [3] ? _01508_ : _01501_;
  assign _01510_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [0] : \MSYNC_1r1w.synth.nz.mem[432] [0];
  assign _01511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [0] : \MSYNC_1r1w.synth.nz.mem[434] [0];
  assign _01512_ = \bapg_rd.w_ptr_r [1] ? _01511_ : _01510_;
  assign _01513_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [0] : \MSYNC_1r1w.synth.nz.mem[436] [0];
  assign _01514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [0] : \MSYNC_1r1w.synth.nz.mem[438] [0];
  assign _01515_ = \bapg_rd.w_ptr_r [1] ? _01514_ : _01513_;
  assign _01516_ = \bapg_rd.w_ptr_r [2] ? _01515_ : _01512_;
  assign _01517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [0] : \MSYNC_1r1w.synth.nz.mem[440] [0];
  assign _01518_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [0] : \MSYNC_1r1w.synth.nz.mem[442] [0];
  assign _01519_ = \bapg_rd.w_ptr_r [1] ? _01518_ : _01517_;
  assign _01520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [0] : \MSYNC_1r1w.synth.nz.mem[444] [0];
  assign _01521_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [0] : \MSYNC_1r1w.synth.nz.mem[446] [0];
  assign _01522_ = \bapg_rd.w_ptr_r [1] ? _01521_ : _01520_;
  assign _01523_ = \bapg_rd.w_ptr_r [2] ? _01522_ : _01519_;
  assign _01524_ = \bapg_rd.w_ptr_r [3] ? _01523_ : _01516_;
  assign _01525_ = \bapg_rd.w_ptr_r [4] ? _01524_ : _01509_;
  assign _01526_ = \bapg_rd.w_ptr_r [5] ? _01525_ : _01494_;
  assign _01527_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [0] : \MSYNC_1r1w.synth.nz.mem[448] [0];
  assign _01528_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [0] : \MSYNC_1r1w.synth.nz.mem[450] [0];
  assign _01529_ = \bapg_rd.w_ptr_r [1] ? _01528_ : _01527_;
  assign _01530_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [0] : \MSYNC_1r1w.synth.nz.mem[452] [0];
  assign _01531_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [0] : \MSYNC_1r1w.synth.nz.mem[454] [0];
  assign _01532_ = \bapg_rd.w_ptr_r [1] ? _01531_ : _01530_;
  assign _01533_ = \bapg_rd.w_ptr_r [2] ? _01532_ : _01529_;
  assign _01534_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [0] : \MSYNC_1r1w.synth.nz.mem[456] [0];
  assign _01535_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [0] : \MSYNC_1r1w.synth.nz.mem[458] [0];
  assign _01536_ = \bapg_rd.w_ptr_r [1] ? _01535_ : _01534_;
  assign _01537_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [0] : \MSYNC_1r1w.synth.nz.mem[460] [0];
  assign _01538_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [0] : \MSYNC_1r1w.synth.nz.mem[462] [0];
  assign _01539_ = \bapg_rd.w_ptr_r [1] ? _01538_ : _01537_;
  assign _01540_ = \bapg_rd.w_ptr_r [2] ? _01539_ : _01536_;
  assign _01541_ = \bapg_rd.w_ptr_r [3] ? _01540_ : _01533_;
  assign _01542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [0] : \MSYNC_1r1w.synth.nz.mem[464] [0];
  assign _01543_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [0] : \MSYNC_1r1w.synth.nz.mem[466] [0];
  assign _01544_ = \bapg_rd.w_ptr_r [1] ? _01543_ : _01542_;
  assign _01545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [0] : \MSYNC_1r1w.synth.nz.mem[468] [0];
  assign _01546_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [0] : \MSYNC_1r1w.synth.nz.mem[470] [0];
  assign _01547_ = \bapg_rd.w_ptr_r [1] ? _01546_ : _01545_;
  assign _01548_ = \bapg_rd.w_ptr_r [2] ? _01547_ : _01544_;
  assign _01549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [0] : \MSYNC_1r1w.synth.nz.mem[472] [0];
  assign _01550_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [0] : \MSYNC_1r1w.synth.nz.mem[474] [0];
  assign _01551_ = \bapg_rd.w_ptr_r [1] ? _01550_ : _01549_;
  assign _01552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [0] : \MSYNC_1r1w.synth.nz.mem[476] [0];
  assign _01553_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [0] : \MSYNC_1r1w.synth.nz.mem[478] [0];
  assign _01554_ = \bapg_rd.w_ptr_r [1] ? _01553_ : _01552_;
  assign _01555_ = \bapg_rd.w_ptr_r [2] ? _01554_ : _01551_;
  assign _01556_ = \bapg_rd.w_ptr_r [3] ? _01555_ : _01548_;
  assign _01557_ = \bapg_rd.w_ptr_r [4] ? _01556_ : _01541_;
  assign _01558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [0] : \MSYNC_1r1w.synth.nz.mem[480] [0];
  assign _01559_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [0] : \MSYNC_1r1w.synth.nz.mem[482] [0];
  assign _01560_ = \bapg_rd.w_ptr_r [1] ? _01559_ : _01558_;
  assign _01561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [0] : \MSYNC_1r1w.synth.nz.mem[484] [0];
  assign _01562_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [0] : \MSYNC_1r1w.synth.nz.mem[486] [0];
  assign _01563_ = \bapg_rd.w_ptr_r [1] ? _01562_ : _01561_;
  assign _01564_ = \bapg_rd.w_ptr_r [2] ? _01563_ : _01560_;
  assign _01565_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [0] : \MSYNC_1r1w.synth.nz.mem[488] [0];
  assign _01566_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [0] : \MSYNC_1r1w.synth.nz.mem[490] [0];
  assign _01567_ = \bapg_rd.w_ptr_r [1] ? _01566_ : _01565_;
  assign _01568_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [0] : \MSYNC_1r1w.synth.nz.mem[492] [0];
  assign _01569_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [0] : \MSYNC_1r1w.synth.nz.mem[494] [0];
  assign _01570_ = \bapg_rd.w_ptr_r [1] ? _01569_ : _01568_;
  assign _01571_ = \bapg_rd.w_ptr_r [2] ? _01570_ : _01567_;
  assign _01572_ = \bapg_rd.w_ptr_r [3] ? _01571_ : _01564_;
  assign _01573_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [0] : \MSYNC_1r1w.synth.nz.mem[496] [0];
  assign _01574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [0] : \MSYNC_1r1w.synth.nz.mem[498] [0];
  assign _01575_ = \bapg_rd.w_ptr_r [1] ? _01574_ : _01573_;
  assign _01576_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [0] : \MSYNC_1r1w.synth.nz.mem[500] [0];
  assign _01577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [0] : \MSYNC_1r1w.synth.nz.mem[502] [0];
  assign _01578_ = \bapg_rd.w_ptr_r [1] ? _01577_ : _01576_;
  assign _01579_ = \bapg_rd.w_ptr_r [2] ? _01578_ : _01575_;
  assign _01580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [0] : \MSYNC_1r1w.synth.nz.mem[504] [0];
  assign _01581_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [0] : \MSYNC_1r1w.synth.nz.mem[506] [0];
  assign _01582_ = \bapg_rd.w_ptr_r [1] ? _01581_ : _01580_;
  assign _01583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [0] : \MSYNC_1r1w.synth.nz.mem[508] [0];
  assign _01584_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [0] : \MSYNC_1r1w.synth.nz.mem[510] [0];
  assign _01585_ = \bapg_rd.w_ptr_r [1] ? _01584_ : _01583_;
  assign _01586_ = \bapg_rd.w_ptr_r [2] ? _01585_ : _01582_;
  assign _01587_ = \bapg_rd.w_ptr_r [3] ? _01586_ : _01579_;
  assign _01588_ = \bapg_rd.w_ptr_r [4] ? _01587_ : _01572_;
  assign _01589_ = \bapg_rd.w_ptr_r [5] ? _01588_ : _01557_;
  assign _01590_ = \bapg_rd.w_ptr_r [6] ? _01589_ : _01526_;
  assign _01591_ = \bapg_rd.w_ptr_r [7] ? _01590_ : _01463_;
  assign _01592_ = \bapg_rd.w_ptr_r [8] ? _01591_ : _01336_;
  assign _01593_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [0] : \MSYNC_1r1w.synth.nz.mem[512] [0];
  assign _01594_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [0] : \MSYNC_1r1w.synth.nz.mem[514] [0];
  assign _01595_ = \bapg_rd.w_ptr_r [1] ? _01594_ : _01593_;
  assign _01596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [0] : \MSYNC_1r1w.synth.nz.mem[516] [0];
  assign _01597_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [0] : \MSYNC_1r1w.synth.nz.mem[518] [0];
  assign _01598_ = \bapg_rd.w_ptr_r [1] ? _01597_ : _01596_;
  assign _01599_ = \bapg_rd.w_ptr_r [2] ? _01598_ : _01595_;
  assign _01600_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [0] : \MSYNC_1r1w.synth.nz.mem[520] [0];
  assign _01601_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [0] : \MSYNC_1r1w.synth.nz.mem[522] [0];
  assign _01602_ = \bapg_rd.w_ptr_r [1] ? _01601_ : _01600_;
  assign _01603_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [0] : \MSYNC_1r1w.synth.nz.mem[524] [0];
  assign _01604_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [0] : \MSYNC_1r1w.synth.nz.mem[526] [0];
  assign _01605_ = \bapg_rd.w_ptr_r [1] ? _01604_ : _01603_;
  assign _01606_ = \bapg_rd.w_ptr_r [2] ? _01605_ : _01602_;
  assign _01607_ = \bapg_rd.w_ptr_r [3] ? _01606_ : _01599_;
  assign _01608_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [0] : \MSYNC_1r1w.synth.nz.mem[528] [0];
  assign _01609_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [0] : \MSYNC_1r1w.synth.nz.mem[530] [0];
  assign _01610_ = \bapg_rd.w_ptr_r [1] ? _01609_ : _01608_;
  assign _01611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [0] : \MSYNC_1r1w.synth.nz.mem[532] [0];
  assign _01612_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [0] : \MSYNC_1r1w.synth.nz.mem[534] [0];
  assign _01613_ = \bapg_rd.w_ptr_r [1] ? _01612_ : _01611_;
  assign _01614_ = \bapg_rd.w_ptr_r [2] ? _01613_ : _01610_;
  assign _01615_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [0] : \MSYNC_1r1w.synth.nz.mem[536] [0];
  assign _01616_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [0] : \MSYNC_1r1w.synth.nz.mem[538] [0];
  assign _01617_ = \bapg_rd.w_ptr_r [1] ? _01616_ : _01615_;
  assign _01618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [0] : \MSYNC_1r1w.synth.nz.mem[540] [0];
  assign _01619_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [0] : \MSYNC_1r1w.synth.nz.mem[542] [0];
  assign _01620_ = \bapg_rd.w_ptr_r [1] ? _01619_ : _01618_;
  assign _01621_ = \bapg_rd.w_ptr_r [2] ? _01620_ : _01617_;
  assign _01622_ = \bapg_rd.w_ptr_r [3] ? _01621_ : _01614_;
  assign _01623_ = \bapg_rd.w_ptr_r [4] ? _01622_ : _01607_;
  assign _01624_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [0] : \MSYNC_1r1w.synth.nz.mem[544] [0];
  assign _01625_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [0] : \MSYNC_1r1w.synth.nz.mem[546] [0];
  assign _01626_ = \bapg_rd.w_ptr_r [1] ? _01625_ : _01624_;
  assign _01627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [0] : \MSYNC_1r1w.synth.nz.mem[548] [0];
  assign _01628_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [0] : \MSYNC_1r1w.synth.nz.mem[550] [0];
  assign _01629_ = \bapg_rd.w_ptr_r [1] ? _01628_ : _01627_;
  assign _01630_ = \bapg_rd.w_ptr_r [2] ? _01629_ : _01626_;
  assign _01631_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [0] : \MSYNC_1r1w.synth.nz.mem[552] [0];
  assign _01632_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [0] : \MSYNC_1r1w.synth.nz.mem[554] [0];
  assign _01633_ = \bapg_rd.w_ptr_r [1] ? _01632_ : _01631_;
  assign _01634_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [0] : \MSYNC_1r1w.synth.nz.mem[556] [0];
  assign _01635_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [0] : \MSYNC_1r1w.synth.nz.mem[558] [0];
  assign _01636_ = \bapg_rd.w_ptr_r [1] ? _01635_ : _01634_;
  assign _01637_ = \bapg_rd.w_ptr_r [2] ? _01636_ : _01633_;
  assign _01638_ = \bapg_rd.w_ptr_r [3] ? _01637_ : _01630_;
  assign _01639_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [0] : \MSYNC_1r1w.synth.nz.mem[560] [0];
  assign _01640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [0] : \MSYNC_1r1w.synth.nz.mem[562] [0];
  assign _01641_ = \bapg_rd.w_ptr_r [1] ? _01640_ : _01639_;
  assign _01642_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [0] : \MSYNC_1r1w.synth.nz.mem[564] [0];
  assign _01643_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [0] : \MSYNC_1r1w.synth.nz.mem[566] [0];
  assign _01644_ = \bapg_rd.w_ptr_r [1] ? _01643_ : _01642_;
  assign _01645_ = \bapg_rd.w_ptr_r [2] ? _01644_ : _01641_;
  assign _01646_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [0] : \MSYNC_1r1w.synth.nz.mem[568] [0];
  assign _01647_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [0] : \MSYNC_1r1w.synth.nz.mem[570] [0];
  assign _01648_ = \bapg_rd.w_ptr_r [1] ? _01647_ : _01646_;
  assign _01649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [0] : \MSYNC_1r1w.synth.nz.mem[572] [0];
  assign _01650_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [0] : \MSYNC_1r1w.synth.nz.mem[574] [0];
  assign _01651_ = \bapg_rd.w_ptr_r [1] ? _01650_ : _01649_;
  assign _01652_ = \bapg_rd.w_ptr_r [2] ? _01651_ : _01648_;
  assign _01653_ = \bapg_rd.w_ptr_r [3] ? _01652_ : _01645_;
  assign _01654_ = \bapg_rd.w_ptr_r [4] ? _01653_ : _01638_;
  assign _01655_ = \bapg_rd.w_ptr_r [5] ? _01654_ : _01623_;
  assign _01656_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [0] : \MSYNC_1r1w.synth.nz.mem[576] [0];
  assign _01657_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [0] : \MSYNC_1r1w.synth.nz.mem[578] [0];
  assign _01658_ = \bapg_rd.w_ptr_r [1] ? _01657_ : _01656_;
  assign _01659_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [0] : \MSYNC_1r1w.synth.nz.mem[580] [0];
  assign _01660_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [0] : \MSYNC_1r1w.synth.nz.mem[582] [0];
  assign _01661_ = \bapg_rd.w_ptr_r [1] ? _01660_ : _01659_;
  assign _01662_ = \bapg_rd.w_ptr_r [2] ? _01661_ : _01658_;
  assign _01663_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [0] : \MSYNC_1r1w.synth.nz.mem[584] [0];
  assign _01664_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [0] : \MSYNC_1r1w.synth.nz.mem[586] [0];
  assign _01665_ = \bapg_rd.w_ptr_r [1] ? _01664_ : _01663_;
  assign _01666_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [0] : \MSYNC_1r1w.synth.nz.mem[588] [0];
  assign _01667_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [0] : \MSYNC_1r1w.synth.nz.mem[590] [0];
  assign _01668_ = \bapg_rd.w_ptr_r [1] ? _01667_ : _01666_;
  assign _01669_ = \bapg_rd.w_ptr_r [2] ? _01668_ : _01665_;
  assign _01670_ = \bapg_rd.w_ptr_r [3] ? _01669_ : _01662_;
  assign _01671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [0] : \MSYNC_1r1w.synth.nz.mem[592] [0];
  assign _01672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [0] : \MSYNC_1r1w.synth.nz.mem[594] [0];
  assign _01673_ = \bapg_rd.w_ptr_r [1] ? _01672_ : _01671_;
  assign _01674_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [0] : \MSYNC_1r1w.synth.nz.mem[596] [0];
  assign _01675_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [0] : \MSYNC_1r1w.synth.nz.mem[598] [0];
  assign _01676_ = \bapg_rd.w_ptr_r [1] ? _01675_ : _01674_;
  assign _01677_ = \bapg_rd.w_ptr_r [2] ? _01676_ : _01673_;
  assign _01678_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [0] : \MSYNC_1r1w.synth.nz.mem[600] [0];
  assign _01679_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [0] : \MSYNC_1r1w.synth.nz.mem[602] [0];
  assign _01680_ = \bapg_rd.w_ptr_r [1] ? _01679_ : _01678_;
  assign _01681_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [0] : \MSYNC_1r1w.synth.nz.mem[604] [0];
  assign _01682_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [0] : \MSYNC_1r1w.synth.nz.mem[606] [0];
  assign _01683_ = \bapg_rd.w_ptr_r [1] ? _01682_ : _01681_;
  assign _01684_ = \bapg_rd.w_ptr_r [2] ? _01683_ : _01680_;
  assign _01685_ = \bapg_rd.w_ptr_r [3] ? _01684_ : _01677_;
  assign _01686_ = \bapg_rd.w_ptr_r [4] ? _01685_ : _01670_;
  assign _01687_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [0] : \MSYNC_1r1w.synth.nz.mem[608] [0];
  assign _01688_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [0] : \MSYNC_1r1w.synth.nz.mem[610] [0];
  assign _01689_ = \bapg_rd.w_ptr_r [1] ? _01688_ : _01687_;
  assign _01690_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [0] : \MSYNC_1r1w.synth.nz.mem[612] [0];
  assign _01691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [0] : \MSYNC_1r1w.synth.nz.mem[614] [0];
  assign _01692_ = \bapg_rd.w_ptr_r [1] ? _01691_ : _01690_;
  assign _01693_ = \bapg_rd.w_ptr_r [2] ? _01692_ : _01689_;
  assign _01694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [0] : \MSYNC_1r1w.synth.nz.mem[616] [0];
  assign _01695_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [0] : \MSYNC_1r1w.synth.nz.mem[618] [0];
  assign _01696_ = \bapg_rd.w_ptr_r [1] ? _01695_ : _01694_;
  assign _01697_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [0] : \MSYNC_1r1w.synth.nz.mem[620] [0];
  assign _01698_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [0] : \MSYNC_1r1w.synth.nz.mem[622] [0];
  assign _01699_ = \bapg_rd.w_ptr_r [1] ? _01698_ : _01697_;
  assign _01700_ = \bapg_rd.w_ptr_r [2] ? _01699_ : _01696_;
  assign _01701_ = \bapg_rd.w_ptr_r [3] ? _01700_ : _01693_;
  assign _01702_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [0] : \MSYNC_1r1w.synth.nz.mem[624] [0];
  assign _01703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [0] : \MSYNC_1r1w.synth.nz.mem[626] [0];
  assign _01704_ = \bapg_rd.w_ptr_r [1] ? _01703_ : _01702_;
  assign _01705_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [0] : \MSYNC_1r1w.synth.nz.mem[628] [0];
  assign _01706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [0] : \MSYNC_1r1w.synth.nz.mem[630] [0];
  assign _01707_ = \bapg_rd.w_ptr_r [1] ? _01706_ : _01705_;
  assign _01708_ = \bapg_rd.w_ptr_r [2] ? _01707_ : _01704_;
  assign _01709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [0] : \MSYNC_1r1w.synth.nz.mem[632] [0];
  assign _01710_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [0] : \MSYNC_1r1w.synth.nz.mem[634] [0];
  assign _01711_ = \bapg_rd.w_ptr_r [1] ? _01710_ : _01709_;
  assign _01712_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [0] : \MSYNC_1r1w.synth.nz.mem[636] [0];
  assign _01713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [0] : \MSYNC_1r1w.synth.nz.mem[638] [0];
  assign _01714_ = \bapg_rd.w_ptr_r [1] ? _01713_ : _01712_;
  assign _01715_ = \bapg_rd.w_ptr_r [2] ? _01714_ : _01711_;
  assign _01716_ = \bapg_rd.w_ptr_r [3] ? _01715_ : _01708_;
  assign _01717_ = \bapg_rd.w_ptr_r [4] ? _01716_ : _01701_;
  assign _01718_ = \bapg_rd.w_ptr_r [5] ? _01717_ : _01686_;
  assign _01719_ = \bapg_rd.w_ptr_r [6] ? _01718_ : _01655_;
  assign _01720_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [0] : \MSYNC_1r1w.synth.nz.mem[640] [0];
  assign _01721_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [0] : \MSYNC_1r1w.synth.nz.mem[642] [0];
  assign _01722_ = \bapg_rd.w_ptr_r [1] ? _01721_ : _01720_;
  assign _01723_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [0] : \MSYNC_1r1w.synth.nz.mem[644] [0];
  assign _01724_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [0] : \MSYNC_1r1w.synth.nz.mem[646] [0];
  assign _01725_ = \bapg_rd.w_ptr_r [1] ? _01724_ : _01723_;
  assign _01726_ = \bapg_rd.w_ptr_r [2] ? _01725_ : _01722_;
  assign _01727_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [0] : \MSYNC_1r1w.synth.nz.mem[648] [0];
  assign _01728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [0] : \MSYNC_1r1w.synth.nz.mem[650] [0];
  assign _01729_ = \bapg_rd.w_ptr_r [1] ? _01728_ : _01727_;
  assign _01730_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [0] : \MSYNC_1r1w.synth.nz.mem[652] [0];
  assign _01731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [0] : \MSYNC_1r1w.synth.nz.mem[654] [0];
  assign _01732_ = \bapg_rd.w_ptr_r [1] ? _01731_ : _01730_;
  assign _01733_ = \bapg_rd.w_ptr_r [2] ? _01732_ : _01729_;
  assign _01734_ = \bapg_rd.w_ptr_r [3] ? _01733_ : _01726_;
  assign _01735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [0] : \MSYNC_1r1w.synth.nz.mem[656] [0];
  assign _01736_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [0] : \MSYNC_1r1w.synth.nz.mem[658] [0];
  assign _01737_ = \bapg_rd.w_ptr_r [1] ? _01736_ : _01735_;
  assign _01738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [0] : \MSYNC_1r1w.synth.nz.mem[660] [0];
  assign _01739_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [0] : \MSYNC_1r1w.synth.nz.mem[662] [0];
  assign _01740_ = \bapg_rd.w_ptr_r [1] ? _01739_ : _01738_;
  assign _01741_ = \bapg_rd.w_ptr_r [2] ? _01740_ : _01737_;
  assign _01742_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [0] : \MSYNC_1r1w.synth.nz.mem[664] [0];
  assign _01743_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [0] : \MSYNC_1r1w.synth.nz.mem[666] [0];
  assign _01744_ = \bapg_rd.w_ptr_r [1] ? _01743_ : _01742_;
  assign _01745_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [0] : \MSYNC_1r1w.synth.nz.mem[668] [0];
  assign _01746_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [0] : \MSYNC_1r1w.synth.nz.mem[670] [0];
  assign _01747_ = \bapg_rd.w_ptr_r [1] ? _01746_ : _01745_;
  assign _01748_ = \bapg_rd.w_ptr_r [2] ? _01747_ : _01744_;
  assign _01749_ = \bapg_rd.w_ptr_r [3] ? _01748_ : _01741_;
  assign _01750_ = \bapg_rd.w_ptr_r [4] ? _01749_ : _01734_;
  assign _01751_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [0] : \MSYNC_1r1w.synth.nz.mem[672] [0];
  assign _01752_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [0] : \MSYNC_1r1w.synth.nz.mem[674] [0];
  assign _01753_ = \bapg_rd.w_ptr_r [1] ? _01752_ : _01751_;
  assign _01754_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [0] : \MSYNC_1r1w.synth.nz.mem[676] [0];
  assign _01755_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [0] : \MSYNC_1r1w.synth.nz.mem[678] [0];
  assign _01756_ = \bapg_rd.w_ptr_r [1] ? _01755_ : _01754_;
  assign _01757_ = \bapg_rd.w_ptr_r [2] ? _01756_ : _01753_;
  assign _01758_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [0] : \MSYNC_1r1w.synth.nz.mem[680] [0];
  assign _01759_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [0] : \MSYNC_1r1w.synth.nz.mem[682] [0];
  assign _01760_ = \bapg_rd.w_ptr_r [1] ? _01759_ : _01758_;
  assign _01761_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [0] : \MSYNC_1r1w.synth.nz.mem[684] [0];
  assign _01762_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [0] : \MSYNC_1r1w.synth.nz.mem[686] [0];
  assign _01763_ = \bapg_rd.w_ptr_r [1] ? _01762_ : _01761_;
  assign _01764_ = \bapg_rd.w_ptr_r [2] ? _01763_ : _01760_;
  assign _01765_ = \bapg_rd.w_ptr_r [3] ? _01764_ : _01757_;
  assign _01766_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [0] : \MSYNC_1r1w.synth.nz.mem[688] [0];
  assign _01767_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [0] : \MSYNC_1r1w.synth.nz.mem[690] [0];
  assign _01768_ = \bapg_rd.w_ptr_r [1] ? _01767_ : _01766_;
  assign _01769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [0] : \MSYNC_1r1w.synth.nz.mem[692] [0];
  assign _01770_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [0] : \MSYNC_1r1w.synth.nz.mem[694] [0];
  assign _01771_ = \bapg_rd.w_ptr_r [1] ? _01770_ : _01769_;
  assign _01772_ = \bapg_rd.w_ptr_r [2] ? _01771_ : _01768_;
  assign _01773_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [0] : \MSYNC_1r1w.synth.nz.mem[696] [0];
  assign _01774_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [0] : \MSYNC_1r1w.synth.nz.mem[698] [0];
  assign _01775_ = \bapg_rd.w_ptr_r [1] ? _01774_ : _01773_;
  assign _01776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [0] : \MSYNC_1r1w.synth.nz.mem[700] [0];
  assign _01777_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [0] : \MSYNC_1r1w.synth.nz.mem[702] [0];
  assign _01778_ = \bapg_rd.w_ptr_r [1] ? _01777_ : _01776_;
  assign _01779_ = \bapg_rd.w_ptr_r [2] ? _01778_ : _01775_;
  assign _01780_ = \bapg_rd.w_ptr_r [3] ? _01779_ : _01772_;
  assign _01781_ = \bapg_rd.w_ptr_r [4] ? _01780_ : _01765_;
  assign _01782_ = \bapg_rd.w_ptr_r [5] ? _01781_ : _01750_;
  assign _01783_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [0] : \MSYNC_1r1w.synth.nz.mem[704] [0];
  assign _01784_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [0] : \MSYNC_1r1w.synth.nz.mem[706] [0];
  assign _01785_ = \bapg_rd.w_ptr_r [1] ? _01784_ : _01783_;
  assign _01786_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [0] : \MSYNC_1r1w.synth.nz.mem[708] [0];
  assign _01787_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [0] : \MSYNC_1r1w.synth.nz.mem[710] [0];
  assign _01788_ = \bapg_rd.w_ptr_r [1] ? _01787_ : _01786_;
  assign _01789_ = \bapg_rd.w_ptr_r [2] ? _01788_ : _01785_;
  assign _01790_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [0] : \MSYNC_1r1w.synth.nz.mem[712] [0];
  assign _01791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [0] : \MSYNC_1r1w.synth.nz.mem[714] [0];
  assign _01792_ = \bapg_rd.w_ptr_r [1] ? _01791_ : _01790_;
  assign _01793_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [0] : \MSYNC_1r1w.synth.nz.mem[716] [0];
  assign _01794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [0] : \MSYNC_1r1w.synth.nz.mem[718] [0];
  assign _01795_ = \bapg_rd.w_ptr_r [1] ? _01794_ : _01793_;
  assign _01796_ = \bapg_rd.w_ptr_r [2] ? _01795_ : _01792_;
  assign _01797_ = \bapg_rd.w_ptr_r [3] ? _01796_ : _01789_;
  assign _01798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [0] : \MSYNC_1r1w.synth.nz.mem[720] [0];
  assign _01799_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [0] : \MSYNC_1r1w.synth.nz.mem[722] [0];
  assign _01800_ = \bapg_rd.w_ptr_r [1] ? _01799_ : _01798_;
  assign _01801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [0] : \MSYNC_1r1w.synth.nz.mem[724] [0];
  assign _01802_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [0] : \MSYNC_1r1w.synth.nz.mem[726] [0];
  assign _01803_ = \bapg_rd.w_ptr_r [1] ? _01802_ : _01801_;
  assign _01804_ = \bapg_rd.w_ptr_r [2] ? _01803_ : _01800_;
  assign _01805_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [0] : \MSYNC_1r1w.synth.nz.mem[728] [0];
  assign _01806_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [0] : \MSYNC_1r1w.synth.nz.mem[730] [0];
  assign _01807_ = \bapg_rd.w_ptr_r [1] ? _01806_ : _01805_;
  assign _01808_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [0] : \MSYNC_1r1w.synth.nz.mem[732] [0];
  assign _01809_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [0] : \MSYNC_1r1w.synth.nz.mem[734] [0];
  assign _01810_ = \bapg_rd.w_ptr_r [1] ? _01809_ : _01808_;
  assign _01811_ = \bapg_rd.w_ptr_r [2] ? _01810_ : _01807_;
  assign _01812_ = \bapg_rd.w_ptr_r [3] ? _01811_ : _01804_;
  assign _01813_ = \bapg_rd.w_ptr_r [4] ? _01812_ : _01797_;
  assign _01814_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [0] : \MSYNC_1r1w.synth.nz.mem[736] [0];
  assign _01815_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [0] : \MSYNC_1r1w.synth.nz.mem[738] [0];
  assign _01816_ = \bapg_rd.w_ptr_r [1] ? _01815_ : _01814_;
  assign _01817_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [0] : \MSYNC_1r1w.synth.nz.mem[740] [0];
  assign _01818_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [0] : \MSYNC_1r1w.synth.nz.mem[742] [0];
  assign _01819_ = \bapg_rd.w_ptr_r [1] ? _01818_ : _01817_;
  assign _01820_ = \bapg_rd.w_ptr_r [2] ? _01819_ : _01816_;
  assign _01821_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [0] : \MSYNC_1r1w.synth.nz.mem[744] [0];
  assign _01822_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [0] : \MSYNC_1r1w.synth.nz.mem[746] [0];
  assign _01823_ = \bapg_rd.w_ptr_r [1] ? _01822_ : _01821_;
  assign _01824_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [0] : \MSYNC_1r1w.synth.nz.mem[748] [0];
  assign _01825_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [0] : \MSYNC_1r1w.synth.nz.mem[750] [0];
  assign _01826_ = \bapg_rd.w_ptr_r [1] ? _01825_ : _01824_;
  assign _01827_ = \bapg_rd.w_ptr_r [2] ? _01826_ : _01823_;
  assign _01828_ = \bapg_rd.w_ptr_r [3] ? _01827_ : _01820_;
  assign _01829_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [0] : \MSYNC_1r1w.synth.nz.mem[752] [0];
  assign _01830_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [0] : \MSYNC_1r1w.synth.nz.mem[754] [0];
  assign _01831_ = \bapg_rd.w_ptr_r [1] ? _01830_ : _01829_;
  assign _01832_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [0] : \MSYNC_1r1w.synth.nz.mem[756] [0];
  assign _01833_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [0] : \MSYNC_1r1w.synth.nz.mem[758] [0];
  assign _01834_ = \bapg_rd.w_ptr_r [1] ? _01833_ : _01832_;
  assign _01835_ = \bapg_rd.w_ptr_r [2] ? _01834_ : _01831_;
  assign _01836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [0] : \MSYNC_1r1w.synth.nz.mem[760] [0];
  assign _01837_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [0] : \MSYNC_1r1w.synth.nz.mem[762] [0];
  assign _01838_ = \bapg_rd.w_ptr_r [1] ? _01837_ : _01836_;
  assign _01839_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [0] : \MSYNC_1r1w.synth.nz.mem[764] [0];
  assign _01840_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [0] : \MSYNC_1r1w.synth.nz.mem[766] [0];
  assign _01841_ = \bapg_rd.w_ptr_r [1] ? _01840_ : _01839_;
  assign _01842_ = \bapg_rd.w_ptr_r [2] ? _01841_ : _01838_;
  assign _01843_ = \bapg_rd.w_ptr_r [3] ? _01842_ : _01835_;
  assign _01844_ = \bapg_rd.w_ptr_r [4] ? _01843_ : _01828_;
  assign _01845_ = \bapg_rd.w_ptr_r [5] ? _01844_ : _01813_;
  assign _01846_ = \bapg_rd.w_ptr_r [6] ? _01845_ : _01782_;
  assign _01847_ = \bapg_rd.w_ptr_r [7] ? _01846_ : _01719_;
  assign _01848_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [0] : \MSYNC_1r1w.synth.nz.mem[768] [0];
  assign _01849_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [0] : \MSYNC_1r1w.synth.nz.mem[770] [0];
  assign _01850_ = \bapg_rd.w_ptr_r [1] ? _01849_ : _01848_;
  assign _01851_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [0] : \MSYNC_1r1w.synth.nz.mem[772] [0];
  assign _01852_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [0] : \MSYNC_1r1w.synth.nz.mem[774] [0];
  assign _01853_ = \bapg_rd.w_ptr_r [1] ? _01852_ : _01851_;
  assign _01854_ = \bapg_rd.w_ptr_r [2] ? _01853_ : _01850_;
  assign _01855_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [0] : \MSYNC_1r1w.synth.nz.mem[776] [0];
  assign _01856_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [0] : \MSYNC_1r1w.synth.nz.mem[778] [0];
  assign _01857_ = \bapg_rd.w_ptr_r [1] ? _01856_ : _01855_;
  assign _01858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [0] : \MSYNC_1r1w.synth.nz.mem[780] [0];
  assign _01859_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [0] : \MSYNC_1r1w.synth.nz.mem[782] [0];
  assign _01860_ = \bapg_rd.w_ptr_r [1] ? _01859_ : _01858_;
  assign _01861_ = \bapg_rd.w_ptr_r [2] ? _01860_ : _01857_;
  assign _01862_ = \bapg_rd.w_ptr_r [3] ? _01861_ : _01854_;
  assign _01863_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [0] : \MSYNC_1r1w.synth.nz.mem[784] [0];
  assign _01864_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [0] : \MSYNC_1r1w.synth.nz.mem[786] [0];
  assign _01865_ = \bapg_rd.w_ptr_r [1] ? _01864_ : _01863_;
  assign _01866_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [0] : \MSYNC_1r1w.synth.nz.mem[788] [0];
  assign _01867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [0] : \MSYNC_1r1w.synth.nz.mem[790] [0];
  assign _01868_ = \bapg_rd.w_ptr_r [1] ? _01867_ : _01866_;
  assign _01869_ = \bapg_rd.w_ptr_r [2] ? _01868_ : _01865_;
  assign _01870_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [0] : \MSYNC_1r1w.synth.nz.mem[792] [0];
  assign _01871_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [0] : \MSYNC_1r1w.synth.nz.mem[794] [0];
  assign _01872_ = \bapg_rd.w_ptr_r [1] ? _01871_ : _01870_;
  assign _01873_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [0] : \MSYNC_1r1w.synth.nz.mem[796] [0];
  assign _01874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [0] : \MSYNC_1r1w.synth.nz.mem[798] [0];
  assign _01875_ = \bapg_rd.w_ptr_r [1] ? _01874_ : _01873_;
  assign _01876_ = \bapg_rd.w_ptr_r [2] ? _01875_ : _01872_;
  assign _01877_ = \bapg_rd.w_ptr_r [3] ? _01876_ : _01869_;
  assign _01878_ = \bapg_rd.w_ptr_r [4] ? _01877_ : _01862_;
  assign _01879_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [0] : \MSYNC_1r1w.synth.nz.mem[800] [0];
  assign _01880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [0] : \MSYNC_1r1w.synth.nz.mem[802] [0];
  assign _01881_ = \bapg_rd.w_ptr_r [1] ? _01880_ : _01879_;
  assign _01882_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [0] : \MSYNC_1r1w.synth.nz.mem[804] [0];
  assign _01883_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [0] : \MSYNC_1r1w.synth.nz.mem[806] [0];
  assign _01884_ = \bapg_rd.w_ptr_r [1] ? _01883_ : _01882_;
  assign _01885_ = \bapg_rd.w_ptr_r [2] ? _01884_ : _01881_;
  assign _01886_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [0] : \MSYNC_1r1w.synth.nz.mem[808] [0];
  assign _01887_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [0] : \MSYNC_1r1w.synth.nz.mem[810] [0];
  assign _01888_ = \bapg_rd.w_ptr_r [1] ? _01887_ : _01886_;
  assign _01889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [0] : \MSYNC_1r1w.synth.nz.mem[812] [0];
  assign _01890_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [0] : \MSYNC_1r1w.synth.nz.mem[814] [0];
  assign _01891_ = \bapg_rd.w_ptr_r [1] ? _01890_ : _01889_;
  assign _01892_ = \bapg_rd.w_ptr_r [2] ? _01891_ : _01888_;
  assign _01893_ = \bapg_rd.w_ptr_r [3] ? _01892_ : _01885_;
  assign _01894_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [0] : \MSYNC_1r1w.synth.nz.mem[816] [0];
  assign _01895_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [0] : \MSYNC_1r1w.synth.nz.mem[818] [0];
  assign _01896_ = \bapg_rd.w_ptr_r [1] ? _01895_ : _01894_;
  assign _01897_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [0] : \MSYNC_1r1w.synth.nz.mem[820] [0];
  assign _01898_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [0] : \MSYNC_1r1w.synth.nz.mem[822] [0];
  assign _01899_ = \bapg_rd.w_ptr_r [1] ? _01898_ : _01897_;
  assign _01900_ = \bapg_rd.w_ptr_r [2] ? _01899_ : _01896_;
  assign _01901_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [0] : \MSYNC_1r1w.synth.nz.mem[824] [0];
  assign _01902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [0] : \MSYNC_1r1w.synth.nz.mem[826] [0];
  assign _01903_ = \bapg_rd.w_ptr_r [1] ? _01902_ : _01901_;
  assign _01904_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [0] : \MSYNC_1r1w.synth.nz.mem[828] [0];
  assign _01905_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [0] : \MSYNC_1r1w.synth.nz.mem[830] [0];
  assign _01906_ = \bapg_rd.w_ptr_r [1] ? _01905_ : _01904_;
  assign _01907_ = \bapg_rd.w_ptr_r [2] ? _01906_ : _01903_;
  assign _01908_ = \bapg_rd.w_ptr_r [3] ? _01907_ : _01900_;
  assign _01909_ = \bapg_rd.w_ptr_r [4] ? _01908_ : _01893_;
  assign _01910_ = \bapg_rd.w_ptr_r [5] ? _01909_ : _01878_;
  assign _01911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [0] : \MSYNC_1r1w.synth.nz.mem[832] [0];
  assign _01912_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [0] : \MSYNC_1r1w.synth.nz.mem[834] [0];
  assign _01913_ = \bapg_rd.w_ptr_r [1] ? _01912_ : _01911_;
  assign _01914_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [0] : \MSYNC_1r1w.synth.nz.mem[836] [0];
  assign _01915_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [0] : \MSYNC_1r1w.synth.nz.mem[838] [0];
  assign _01916_ = \bapg_rd.w_ptr_r [1] ? _01915_ : _01914_;
  assign _01917_ = \bapg_rd.w_ptr_r [2] ? _01916_ : _01913_;
  assign _01918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [0] : \MSYNC_1r1w.synth.nz.mem[840] [0];
  assign _01919_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [0] : \MSYNC_1r1w.synth.nz.mem[842] [0];
  assign _01920_ = \bapg_rd.w_ptr_r [1] ? _01919_ : _01918_;
  assign _01921_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [0] : \MSYNC_1r1w.synth.nz.mem[844] [0];
  assign _01922_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [0] : \MSYNC_1r1w.synth.nz.mem[846] [0];
  assign _01923_ = \bapg_rd.w_ptr_r [1] ? _01922_ : _01921_;
  assign _01924_ = \bapg_rd.w_ptr_r [2] ? _01923_ : _01920_;
  assign _01925_ = \bapg_rd.w_ptr_r [3] ? _01924_ : _01917_;
  assign _01926_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [0] : \MSYNC_1r1w.synth.nz.mem[848] [0];
  assign _01927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [0] : \MSYNC_1r1w.synth.nz.mem[850] [0];
  assign _01928_ = \bapg_rd.w_ptr_r [1] ? _01927_ : _01926_;
  assign _01929_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [0] : \MSYNC_1r1w.synth.nz.mem[852] [0];
  assign _01930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [0] : \MSYNC_1r1w.synth.nz.mem[854] [0];
  assign _01931_ = \bapg_rd.w_ptr_r [1] ? _01930_ : _01929_;
  assign _01932_ = \bapg_rd.w_ptr_r [2] ? _01931_ : _01928_;
  assign _01933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [0] : \MSYNC_1r1w.synth.nz.mem[856] [0];
  assign _01934_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [0] : \MSYNC_1r1w.synth.nz.mem[858] [0];
  assign _01935_ = \bapg_rd.w_ptr_r [1] ? _01934_ : _01933_;
  assign _01936_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [0] : \MSYNC_1r1w.synth.nz.mem[860] [0];
  assign _01937_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [0] : \MSYNC_1r1w.synth.nz.mem[862] [0];
  assign _01938_ = \bapg_rd.w_ptr_r [1] ? _01937_ : _01936_;
  assign _01939_ = \bapg_rd.w_ptr_r [2] ? _01938_ : _01935_;
  assign _01940_ = \bapg_rd.w_ptr_r [3] ? _01939_ : _01932_;
  assign _01941_ = \bapg_rd.w_ptr_r [4] ? _01940_ : _01925_;
  assign _01942_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [0] : \MSYNC_1r1w.synth.nz.mem[864] [0];
  assign _01943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [0] : \MSYNC_1r1w.synth.nz.mem[866] [0];
  assign _01944_ = \bapg_rd.w_ptr_r [1] ? _01943_ : _01942_;
  assign _01945_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [0] : \MSYNC_1r1w.synth.nz.mem[868] [0];
  assign _01946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [0] : \MSYNC_1r1w.synth.nz.mem[870] [0];
  assign _01947_ = \bapg_rd.w_ptr_r [1] ? _01946_ : _01945_;
  assign _01948_ = \bapg_rd.w_ptr_r [2] ? _01947_ : _01944_;
  assign _01949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [0] : \MSYNC_1r1w.synth.nz.mem[872] [0];
  assign _01950_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [0] : \MSYNC_1r1w.synth.nz.mem[874] [0];
  assign _01951_ = \bapg_rd.w_ptr_r [1] ? _01950_ : _01949_;
  assign _01952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [0] : \MSYNC_1r1w.synth.nz.mem[876] [0];
  assign _01953_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [0] : \MSYNC_1r1w.synth.nz.mem[878] [0];
  assign _01954_ = \bapg_rd.w_ptr_r [1] ? _01953_ : _01952_;
  assign _01955_ = \bapg_rd.w_ptr_r [2] ? _01954_ : _01951_;
  assign _01956_ = \bapg_rd.w_ptr_r [3] ? _01955_ : _01948_;
  assign _01957_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [0] : \MSYNC_1r1w.synth.nz.mem[880] [0];
  assign _01958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [0] : \MSYNC_1r1w.synth.nz.mem[882] [0];
  assign _01959_ = \bapg_rd.w_ptr_r [1] ? _01958_ : _01957_;
  assign _01960_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [0] : \MSYNC_1r1w.synth.nz.mem[884] [0];
  assign _01961_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [0] : \MSYNC_1r1w.synth.nz.mem[886] [0];
  assign _01962_ = \bapg_rd.w_ptr_r [1] ? _01961_ : _01960_;
  assign _01963_ = \bapg_rd.w_ptr_r [2] ? _01962_ : _01959_;
  assign _01964_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [0] : \MSYNC_1r1w.synth.nz.mem[888] [0];
  assign _01965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [0] : \MSYNC_1r1w.synth.nz.mem[890] [0];
  assign _01966_ = \bapg_rd.w_ptr_r [1] ? _01965_ : _01964_;
  assign _01967_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [0] : \MSYNC_1r1w.synth.nz.mem[892] [0];
  assign _01968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [0] : \MSYNC_1r1w.synth.nz.mem[894] [0];
  assign _01969_ = \bapg_rd.w_ptr_r [1] ? _01968_ : _01967_;
  assign _01970_ = \bapg_rd.w_ptr_r [2] ? _01969_ : _01966_;
  assign _01971_ = \bapg_rd.w_ptr_r [3] ? _01970_ : _01963_;
  assign _01972_ = \bapg_rd.w_ptr_r [4] ? _01971_ : _01956_;
  assign _01973_ = \bapg_rd.w_ptr_r [5] ? _01972_ : _01941_;
  assign _01974_ = \bapg_rd.w_ptr_r [6] ? _01973_ : _01910_;
  assign _01975_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [0] : \MSYNC_1r1w.synth.nz.mem[896] [0];
  assign _01976_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [0] : \MSYNC_1r1w.synth.nz.mem[898] [0];
  assign _01977_ = \bapg_rd.w_ptr_r [1] ? _01976_ : _01975_;
  assign _01978_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [0] : \MSYNC_1r1w.synth.nz.mem[900] [0];
  assign _01979_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [0] : \MSYNC_1r1w.synth.nz.mem[902] [0];
  assign _01980_ = \bapg_rd.w_ptr_r [1] ? _01979_ : _01978_;
  assign _01981_ = \bapg_rd.w_ptr_r [2] ? _01980_ : _01977_;
  assign _01982_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [0] : \MSYNC_1r1w.synth.nz.mem[904] [0];
  assign _01983_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [0] : \MSYNC_1r1w.synth.nz.mem[906] [0];
  assign _01984_ = \bapg_rd.w_ptr_r [1] ? _01983_ : _01982_;
  assign _01985_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [0] : \MSYNC_1r1w.synth.nz.mem[908] [0];
  assign _01986_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [0] : \MSYNC_1r1w.synth.nz.mem[910] [0];
  assign _01987_ = \bapg_rd.w_ptr_r [1] ? _01986_ : _01985_;
  assign _01988_ = \bapg_rd.w_ptr_r [2] ? _01987_ : _01984_;
  assign _01989_ = \bapg_rd.w_ptr_r [3] ? _01988_ : _01981_;
  assign _01990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [0] : \MSYNC_1r1w.synth.nz.mem[912] [0];
  assign _01991_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [0] : \MSYNC_1r1w.synth.nz.mem[914] [0];
  assign _01992_ = \bapg_rd.w_ptr_r [1] ? _01991_ : _01990_;
  assign _01993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [0] : \MSYNC_1r1w.synth.nz.mem[916] [0];
  assign _01994_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [0] : \MSYNC_1r1w.synth.nz.mem[918] [0];
  assign _01995_ = \bapg_rd.w_ptr_r [1] ? _01994_ : _01993_;
  assign _01996_ = \bapg_rd.w_ptr_r [2] ? _01995_ : _01992_;
  assign _01997_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [0] : \MSYNC_1r1w.synth.nz.mem[920] [0];
  assign _01998_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [0] : \MSYNC_1r1w.synth.nz.mem[922] [0];
  assign _01999_ = \bapg_rd.w_ptr_r [1] ? _01998_ : _01997_;
  assign _02000_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [0] : \MSYNC_1r1w.synth.nz.mem[924] [0];
  assign _02001_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [0] : \MSYNC_1r1w.synth.nz.mem[926] [0];
  assign _02002_ = \bapg_rd.w_ptr_r [1] ? _02001_ : _02000_;
  assign _02003_ = \bapg_rd.w_ptr_r [2] ? _02002_ : _01999_;
  assign _02004_ = \bapg_rd.w_ptr_r [3] ? _02003_ : _01996_;
  assign _02005_ = \bapg_rd.w_ptr_r [4] ? _02004_ : _01989_;
  assign _02006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [0] : \MSYNC_1r1w.synth.nz.mem[928] [0];
  assign _02007_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [0] : \MSYNC_1r1w.synth.nz.mem[930] [0];
  assign _02008_ = \bapg_rd.w_ptr_r [1] ? _02007_ : _02006_;
  assign _02009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [0] : \MSYNC_1r1w.synth.nz.mem[932] [0];
  assign _02010_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [0] : \MSYNC_1r1w.synth.nz.mem[934] [0];
  assign _02011_ = \bapg_rd.w_ptr_r [1] ? _02010_ : _02009_;
  assign _02012_ = \bapg_rd.w_ptr_r [2] ? _02011_ : _02008_;
  assign _02013_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [0] : \MSYNC_1r1w.synth.nz.mem[936] [0];
  assign _02014_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [0] : \MSYNC_1r1w.synth.nz.mem[938] [0];
  assign _02015_ = \bapg_rd.w_ptr_r [1] ? _02014_ : _02013_;
  assign _02016_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [0] : \MSYNC_1r1w.synth.nz.mem[940] [0];
  assign _02017_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [0] : \MSYNC_1r1w.synth.nz.mem[942] [0];
  assign _02018_ = \bapg_rd.w_ptr_r [1] ? _02017_ : _02016_;
  assign _02019_ = \bapg_rd.w_ptr_r [2] ? _02018_ : _02015_;
  assign _02020_ = \bapg_rd.w_ptr_r [3] ? _02019_ : _02012_;
  assign _02021_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [0] : \MSYNC_1r1w.synth.nz.mem[944] [0];
  assign _02022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [0] : \MSYNC_1r1w.synth.nz.mem[946] [0];
  assign _02023_ = \bapg_rd.w_ptr_r [1] ? _02022_ : _02021_;
  assign _02024_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [0] : \MSYNC_1r1w.synth.nz.mem[948] [0];
  assign _02025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [0] : \MSYNC_1r1w.synth.nz.mem[950] [0];
  assign _02026_ = \bapg_rd.w_ptr_r [1] ? _02025_ : _02024_;
  assign _02027_ = \bapg_rd.w_ptr_r [2] ? _02026_ : _02023_;
  assign _02028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [0] : \MSYNC_1r1w.synth.nz.mem[952] [0];
  assign _02029_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [0] : \MSYNC_1r1w.synth.nz.mem[954] [0];
  assign _02030_ = \bapg_rd.w_ptr_r [1] ? _02029_ : _02028_;
  assign _02031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [0] : \MSYNC_1r1w.synth.nz.mem[956] [0];
  assign _02032_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [0] : \MSYNC_1r1w.synth.nz.mem[958] [0];
  assign _02033_ = \bapg_rd.w_ptr_r [1] ? _02032_ : _02031_;
  assign _02034_ = \bapg_rd.w_ptr_r [2] ? _02033_ : _02030_;
  assign _02035_ = \bapg_rd.w_ptr_r [3] ? _02034_ : _02027_;
  assign _02036_ = \bapg_rd.w_ptr_r [4] ? _02035_ : _02020_;
  assign _02037_ = \bapg_rd.w_ptr_r [5] ? _02036_ : _02005_;
  assign _02038_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [0] : \MSYNC_1r1w.synth.nz.mem[960] [0];
  assign _02039_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [0] : \MSYNC_1r1w.synth.nz.mem[962] [0];
  assign _02040_ = \bapg_rd.w_ptr_r [1] ? _02039_ : _02038_;
  assign _02041_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [0] : \MSYNC_1r1w.synth.nz.mem[964] [0];
  assign _02042_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [0] : \MSYNC_1r1w.synth.nz.mem[966] [0];
  assign _02043_ = \bapg_rd.w_ptr_r [1] ? _02042_ : _02041_;
  assign _02044_ = \bapg_rd.w_ptr_r [2] ? _02043_ : _02040_;
  assign _02045_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [0] : \MSYNC_1r1w.synth.nz.mem[968] [0];
  assign _02046_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [0] : \MSYNC_1r1w.synth.nz.mem[970] [0];
  assign _02047_ = \bapg_rd.w_ptr_r [1] ? _02046_ : _02045_;
  assign _02048_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [0] : \MSYNC_1r1w.synth.nz.mem[972] [0];
  assign _02049_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [0] : \MSYNC_1r1w.synth.nz.mem[974] [0];
  assign _02050_ = \bapg_rd.w_ptr_r [1] ? _02049_ : _02048_;
  assign _02051_ = \bapg_rd.w_ptr_r [2] ? _02050_ : _02047_;
  assign _02052_ = \bapg_rd.w_ptr_r [3] ? _02051_ : _02044_;
  assign _02053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [0] : \MSYNC_1r1w.synth.nz.mem[976] [0];
  assign _02054_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [0] : \MSYNC_1r1w.synth.nz.mem[978] [0];
  assign _02055_ = \bapg_rd.w_ptr_r [1] ? _02054_ : _02053_;
  assign _02056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [0] : \MSYNC_1r1w.synth.nz.mem[980] [0];
  assign _02057_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [0] : \MSYNC_1r1w.synth.nz.mem[982] [0];
  assign _02058_ = \bapg_rd.w_ptr_r [1] ? _02057_ : _02056_;
  assign _02059_ = \bapg_rd.w_ptr_r [2] ? _02058_ : _02055_;
  assign _02060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [0] : \MSYNC_1r1w.synth.nz.mem[984] [0];
  assign _02061_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [0] : \MSYNC_1r1w.synth.nz.mem[986] [0];
  assign _02062_ = \bapg_rd.w_ptr_r [1] ? _02061_ : _02060_;
  assign _02063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [0] : \MSYNC_1r1w.synth.nz.mem[988] [0];
  assign _02064_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [0] : \MSYNC_1r1w.synth.nz.mem[990] [0];
  assign _02065_ = \bapg_rd.w_ptr_r [1] ? _02064_ : _02063_;
  assign _02066_ = \bapg_rd.w_ptr_r [2] ? _02065_ : _02062_;
  assign _02067_ = \bapg_rd.w_ptr_r [3] ? _02066_ : _02059_;
  assign _02068_ = \bapg_rd.w_ptr_r [4] ? _02067_ : _02052_;
  assign _02069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [0] : \MSYNC_1r1w.synth.nz.mem[992] [0];
  assign _02070_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [0] : \MSYNC_1r1w.synth.nz.mem[994] [0];
  assign _02071_ = \bapg_rd.w_ptr_r [1] ? _02070_ : _02069_;
  assign _02072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [0] : \MSYNC_1r1w.synth.nz.mem[996] [0];
  assign _02073_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [0] : \MSYNC_1r1w.synth.nz.mem[998] [0];
  assign _02074_ = \bapg_rd.w_ptr_r [1] ? _02073_ : _02072_;
  assign _02075_ = \bapg_rd.w_ptr_r [2] ? _02074_ : _02071_;
  assign _02076_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [0] : \MSYNC_1r1w.synth.nz.mem[1000] [0];
  assign _02077_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [0] : \MSYNC_1r1w.synth.nz.mem[1002] [0];
  assign _02078_ = \bapg_rd.w_ptr_r [1] ? _02077_ : _02076_;
  assign _02079_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [0] : \MSYNC_1r1w.synth.nz.mem[1004] [0];
  assign _02080_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [0] : \MSYNC_1r1w.synth.nz.mem[1006] [0];
  assign _02081_ = \bapg_rd.w_ptr_r [1] ? _02080_ : _02079_;
  assign _02082_ = \bapg_rd.w_ptr_r [2] ? _02081_ : _02078_;
  assign _02083_ = \bapg_rd.w_ptr_r [3] ? _02082_ : _02075_;
  assign _02084_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [0] : \MSYNC_1r1w.synth.nz.mem[1008] [0];
  assign _02085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [0] : \MSYNC_1r1w.synth.nz.mem[1010] [0];
  assign _02086_ = \bapg_rd.w_ptr_r [1] ? _02085_ : _02084_;
  assign _02087_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [0] : \MSYNC_1r1w.synth.nz.mem[1012] [0];
  assign _02088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [0] : \MSYNC_1r1w.synth.nz.mem[1014] [0];
  assign _02089_ = \bapg_rd.w_ptr_r [1] ? _02088_ : _02087_;
  assign _02090_ = \bapg_rd.w_ptr_r [2] ? _02089_ : _02086_;
  assign _02091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [0] : \MSYNC_1r1w.synth.nz.mem[1016] [0];
  assign _02092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [0] : \MSYNC_1r1w.synth.nz.mem[1018] [0];
  assign _02093_ = \bapg_rd.w_ptr_r [1] ? _02092_ : _02091_;
  assign _02094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [0] : \MSYNC_1r1w.synth.nz.mem[1020] [0];
  assign _02095_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [0] : \MSYNC_1r1w.synth.nz.mem[1022] [0];
  assign _02096_ = \bapg_rd.w_ptr_r [1] ? _02095_ : _02094_;
  assign _02097_ = \bapg_rd.w_ptr_r [2] ? _02096_ : _02093_;
  assign _02098_ = \bapg_rd.w_ptr_r [3] ? _02097_ : _02090_;
  assign _02099_ = \bapg_rd.w_ptr_r [4] ? _02098_ : _02083_;
  assign _02100_ = \bapg_rd.w_ptr_r [5] ? _02099_ : _02068_;
  assign _02101_ = \bapg_rd.w_ptr_r [6] ? _02100_ : _02037_;
  assign _02102_ = \bapg_rd.w_ptr_r [7] ? _02101_ : _01974_;
  assign _02103_ = \bapg_rd.w_ptr_r [8] ? _02102_ : _01847_;
  assign r_data_o[0] = \bapg_rd.w_ptr_r [9] ? _02103_ : _01592_;
  assign _02104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [1] : \MSYNC_1r1w.synth.nz.mem[0] [1];
  assign _02105_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [1] : \MSYNC_1r1w.synth.nz.mem[2] [1];
  assign _02106_ = \bapg_rd.w_ptr_r [1] ? _02105_ : _02104_;
  assign _02107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [1] : \MSYNC_1r1w.synth.nz.mem[4] [1];
  assign _02108_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [1] : \MSYNC_1r1w.synth.nz.mem[6] [1];
  assign _02109_ = \bapg_rd.w_ptr_r [1] ? _02108_ : _02107_;
  assign _02110_ = \bapg_rd.w_ptr_r [2] ? _02109_ : _02106_;
  assign _02111_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [1] : \MSYNC_1r1w.synth.nz.mem[8] [1];
  assign _02112_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [1] : \MSYNC_1r1w.synth.nz.mem[10] [1];
  assign _02113_ = \bapg_rd.w_ptr_r [1] ? _02112_ : _02111_;
  assign _02114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [1] : \MSYNC_1r1w.synth.nz.mem[12] [1];
  assign _02115_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [1] : \MSYNC_1r1w.synth.nz.mem[14] [1];
  assign _02116_ = \bapg_rd.w_ptr_r [1] ? _02115_ : _02114_;
  assign _02117_ = \bapg_rd.w_ptr_r [2] ? _02116_ : _02113_;
  assign _02118_ = \bapg_rd.w_ptr_r [3] ? _02117_ : _02110_;
  assign _02119_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [1] : \MSYNC_1r1w.synth.nz.mem[16] [1];
  assign _02120_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [1] : \MSYNC_1r1w.synth.nz.mem[18] [1];
  assign _02121_ = \bapg_rd.w_ptr_r [1] ? _02120_ : _02119_;
  assign _02122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [1] : \MSYNC_1r1w.synth.nz.mem[20] [1];
  assign _02123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [1] : \MSYNC_1r1w.synth.nz.mem[22] [1];
  assign _02124_ = \bapg_rd.w_ptr_r [1] ? _02123_ : _02122_;
  assign _02125_ = \bapg_rd.w_ptr_r [2] ? _02124_ : _02121_;
  assign _02126_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [1] : \MSYNC_1r1w.synth.nz.mem[24] [1];
  assign _02127_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [1] : \MSYNC_1r1w.synth.nz.mem[26] [1];
  assign _02128_ = \bapg_rd.w_ptr_r [1] ? _02127_ : _02126_;
  assign _02129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [1] : \MSYNC_1r1w.synth.nz.mem[28] [1];
  assign _02130_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [1] : \MSYNC_1r1w.synth.nz.mem[30] [1];
  assign _02131_ = \bapg_rd.w_ptr_r [1] ? _02130_ : _02129_;
  assign _02132_ = \bapg_rd.w_ptr_r [2] ? _02131_ : _02128_;
  assign _02133_ = \bapg_rd.w_ptr_r [3] ? _02132_ : _02125_;
  assign _02134_ = \bapg_rd.w_ptr_r [4] ? _02133_ : _02118_;
  assign _02135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [1] : \MSYNC_1r1w.synth.nz.mem[32] [1];
  assign _02136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [1] : \MSYNC_1r1w.synth.nz.mem[34] [1];
  assign _02137_ = \bapg_rd.w_ptr_r [1] ? _02136_ : _02135_;
  assign _02138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [1] : \MSYNC_1r1w.synth.nz.mem[36] [1];
  assign _02139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [1] : \MSYNC_1r1w.synth.nz.mem[38] [1];
  assign _02140_ = \bapg_rd.w_ptr_r [1] ? _02139_ : _02138_;
  assign _02141_ = \bapg_rd.w_ptr_r [2] ? _02140_ : _02137_;
  assign _02142_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [1] : \MSYNC_1r1w.synth.nz.mem[40] [1];
  assign _02143_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [1] : \MSYNC_1r1w.synth.nz.mem[42] [1];
  assign _02144_ = \bapg_rd.w_ptr_r [1] ? _02143_ : _02142_;
  assign _02145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [1] : \MSYNC_1r1w.synth.nz.mem[44] [1];
  assign _02146_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [1] : \MSYNC_1r1w.synth.nz.mem[46] [1];
  assign _02147_ = \bapg_rd.w_ptr_r [1] ? _02146_ : _02145_;
  assign _02148_ = \bapg_rd.w_ptr_r [2] ? _02147_ : _02144_;
  assign _02149_ = \bapg_rd.w_ptr_r [3] ? _02148_ : _02141_;
  assign _02150_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [1] : \MSYNC_1r1w.synth.nz.mem[48] [1];
  assign _02151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [1] : \MSYNC_1r1w.synth.nz.mem[50] [1];
  assign _02152_ = \bapg_rd.w_ptr_r [1] ? _02151_ : _02150_;
  assign _02153_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [1] : \MSYNC_1r1w.synth.nz.mem[52] [1];
  assign _02154_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [1] : \MSYNC_1r1w.synth.nz.mem[54] [1];
  assign _02155_ = \bapg_rd.w_ptr_r [1] ? _02154_ : _02153_;
  assign _02156_ = \bapg_rd.w_ptr_r [2] ? _02155_ : _02152_;
  assign _02157_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [1] : \MSYNC_1r1w.synth.nz.mem[56] [1];
  assign _02158_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [1] : \MSYNC_1r1w.synth.nz.mem[58] [1];
  assign _02159_ = \bapg_rd.w_ptr_r [1] ? _02158_ : _02157_;
  assign _02160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [1] : \MSYNC_1r1w.synth.nz.mem[60] [1];
  assign _02161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [1] : \MSYNC_1r1w.synth.nz.mem[62] [1];
  assign _02162_ = \bapg_rd.w_ptr_r [1] ? _02161_ : _02160_;
  assign _02163_ = \bapg_rd.w_ptr_r [2] ? _02162_ : _02159_;
  assign _02164_ = \bapg_rd.w_ptr_r [3] ? _02163_ : _02156_;
  assign _02165_ = \bapg_rd.w_ptr_r [4] ? _02164_ : _02149_;
  assign _02166_ = \bapg_rd.w_ptr_r [5] ? _02165_ : _02134_;
  assign _02167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [1] : \MSYNC_1r1w.synth.nz.mem[64] [1];
  assign _02168_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [1] : \MSYNC_1r1w.synth.nz.mem[66] [1];
  assign _02169_ = \bapg_rd.w_ptr_r [1] ? _02168_ : _02167_;
  assign _02170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [1] : \MSYNC_1r1w.synth.nz.mem[68] [1];
  assign _02171_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [1] : \MSYNC_1r1w.synth.nz.mem[70] [1];
  assign _02172_ = \bapg_rd.w_ptr_r [1] ? _02171_ : _02170_;
  assign _02173_ = \bapg_rd.w_ptr_r [2] ? _02172_ : _02169_;
  assign _02174_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [1] : \MSYNC_1r1w.synth.nz.mem[72] [1];
  assign _02175_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [1] : \MSYNC_1r1w.synth.nz.mem[74] [1];
  assign _02176_ = \bapg_rd.w_ptr_r [1] ? _02175_ : _02174_;
  assign _02177_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [1] : \MSYNC_1r1w.synth.nz.mem[76] [1];
  assign _02178_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [1] : \MSYNC_1r1w.synth.nz.mem[78] [1];
  assign _02179_ = \bapg_rd.w_ptr_r [1] ? _02178_ : _02177_;
  assign _02180_ = \bapg_rd.w_ptr_r [2] ? _02179_ : _02176_;
  assign _02181_ = \bapg_rd.w_ptr_r [3] ? _02180_ : _02173_;
  assign _02182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [1] : \MSYNC_1r1w.synth.nz.mem[80] [1];
  assign _02183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [1] : \MSYNC_1r1w.synth.nz.mem[82] [1];
  assign _02184_ = \bapg_rd.w_ptr_r [1] ? _02183_ : _02182_;
  assign _02185_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [1] : \MSYNC_1r1w.synth.nz.mem[84] [1];
  assign _02186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [1] : \MSYNC_1r1w.synth.nz.mem[86] [1];
  assign _02187_ = \bapg_rd.w_ptr_r [1] ? _02186_ : _02185_;
  assign _02188_ = \bapg_rd.w_ptr_r [2] ? _02187_ : _02184_;
  assign _02189_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [1] : \MSYNC_1r1w.synth.nz.mem[88] [1];
  assign _02190_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [1] : \MSYNC_1r1w.synth.nz.mem[90] [1];
  assign _02191_ = \bapg_rd.w_ptr_r [1] ? _02190_ : _02189_;
  assign _02192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [1] : \MSYNC_1r1w.synth.nz.mem[92] [1];
  assign _02193_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [1] : \MSYNC_1r1w.synth.nz.mem[94] [1];
  assign _02194_ = \bapg_rd.w_ptr_r [1] ? _02193_ : _02192_;
  assign _02195_ = \bapg_rd.w_ptr_r [2] ? _02194_ : _02191_;
  assign _02196_ = \bapg_rd.w_ptr_r [3] ? _02195_ : _02188_;
  assign _02197_ = \bapg_rd.w_ptr_r [4] ? _02196_ : _02181_;
  assign _02198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [1] : \MSYNC_1r1w.synth.nz.mem[96] [1];
  assign _02199_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [1] : \MSYNC_1r1w.synth.nz.mem[98] [1];
  assign _02200_ = \bapg_rd.w_ptr_r [1] ? _02199_ : _02198_;
  assign _02201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [1] : \MSYNC_1r1w.synth.nz.mem[100] [1];
  assign _02202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [1] : \MSYNC_1r1w.synth.nz.mem[102] [1];
  assign _02203_ = \bapg_rd.w_ptr_r [1] ? _02202_ : _02201_;
  assign _02204_ = \bapg_rd.w_ptr_r [2] ? _02203_ : _02200_;
  assign _02205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [1] : \MSYNC_1r1w.synth.nz.mem[104] [1];
  assign _02206_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [1] : \MSYNC_1r1w.synth.nz.mem[106] [1];
  assign _02207_ = \bapg_rd.w_ptr_r [1] ? _02206_ : _02205_;
  assign _02208_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [1] : \MSYNC_1r1w.synth.nz.mem[108] [1];
  assign _02209_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [1] : \MSYNC_1r1w.synth.nz.mem[110] [1];
  assign _02210_ = \bapg_rd.w_ptr_r [1] ? _02209_ : _02208_;
  assign _02211_ = \bapg_rd.w_ptr_r [2] ? _02210_ : _02207_;
  assign _02212_ = \bapg_rd.w_ptr_r [3] ? _02211_ : _02204_;
  assign _02213_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [1] : \MSYNC_1r1w.synth.nz.mem[112] [1];
  assign _02214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [1] : \MSYNC_1r1w.synth.nz.mem[114] [1];
  assign _02215_ = \bapg_rd.w_ptr_r [1] ? _02214_ : _02213_;
  assign _02216_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [1] : \MSYNC_1r1w.synth.nz.mem[116] [1];
  assign _02217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [1] : \MSYNC_1r1w.synth.nz.mem[118] [1];
  assign _02218_ = \bapg_rd.w_ptr_r [1] ? _02217_ : _02216_;
  assign _02219_ = \bapg_rd.w_ptr_r [2] ? _02218_ : _02215_;
  assign _02220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [1] : \MSYNC_1r1w.synth.nz.mem[120] [1];
  assign _02221_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [1] : \MSYNC_1r1w.synth.nz.mem[122] [1];
  assign _02222_ = \bapg_rd.w_ptr_r [1] ? _02221_ : _02220_;
  assign _02223_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [1] : \MSYNC_1r1w.synth.nz.mem[124] [1];
  assign _02224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [1] : \MSYNC_1r1w.synth.nz.mem[126] [1];
  assign _02225_ = \bapg_rd.w_ptr_r [1] ? _02224_ : _02223_;
  assign _02226_ = \bapg_rd.w_ptr_r [2] ? _02225_ : _02222_;
  assign _02227_ = \bapg_rd.w_ptr_r [3] ? _02226_ : _02219_;
  assign _02228_ = \bapg_rd.w_ptr_r [4] ? _02227_ : _02212_;
  assign _02229_ = \bapg_rd.w_ptr_r [5] ? _02228_ : _02197_;
  assign _02230_ = \bapg_rd.w_ptr_r [6] ? _02229_ : _02166_;
  assign _02231_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [1] : \MSYNC_1r1w.synth.nz.mem[128] [1];
  assign _02232_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [1] : \MSYNC_1r1w.synth.nz.mem[130] [1];
  assign _02233_ = \bapg_rd.w_ptr_r [1] ? _02232_ : _02231_;
  assign _02234_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [1] : \MSYNC_1r1w.synth.nz.mem[132] [1];
  assign _02235_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [1] : \MSYNC_1r1w.synth.nz.mem[134] [1];
  assign _02236_ = \bapg_rd.w_ptr_r [1] ? _02235_ : _02234_;
  assign _02237_ = \bapg_rd.w_ptr_r [2] ? _02236_ : _02233_;
  assign _02238_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [1] : \MSYNC_1r1w.synth.nz.mem[136] [1];
  assign _02239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [1] : \MSYNC_1r1w.synth.nz.mem[138] [1];
  assign _02240_ = \bapg_rd.w_ptr_r [1] ? _02239_ : _02238_;
  assign _02241_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [1] : \MSYNC_1r1w.synth.nz.mem[140] [1];
  assign _02242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [1] : \MSYNC_1r1w.synth.nz.mem[142] [1];
  assign _02243_ = \bapg_rd.w_ptr_r [1] ? _02242_ : _02241_;
  assign _02244_ = \bapg_rd.w_ptr_r [2] ? _02243_ : _02240_;
  assign _02245_ = \bapg_rd.w_ptr_r [3] ? _02244_ : _02237_;
  assign _02246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [1] : \MSYNC_1r1w.synth.nz.mem[144] [1];
  assign _02247_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [1] : \MSYNC_1r1w.synth.nz.mem[146] [1];
  assign _02248_ = \bapg_rd.w_ptr_r [1] ? _02247_ : _02246_;
  assign _02249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [1] : \MSYNC_1r1w.synth.nz.mem[148] [1];
  assign _02250_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [1] : \MSYNC_1r1w.synth.nz.mem[150] [1];
  assign _02251_ = \bapg_rd.w_ptr_r [1] ? _02250_ : _02249_;
  assign _02252_ = \bapg_rd.w_ptr_r [2] ? _02251_ : _02248_;
  assign _02253_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [1] : \MSYNC_1r1w.synth.nz.mem[152] [1];
  assign _02254_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [1] : \MSYNC_1r1w.synth.nz.mem[154] [1];
  assign _02255_ = \bapg_rd.w_ptr_r [1] ? _02254_ : _02253_;
  assign _02256_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [1] : \MSYNC_1r1w.synth.nz.mem[156] [1];
  assign _02257_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [1] : \MSYNC_1r1w.synth.nz.mem[158] [1];
  assign _02258_ = \bapg_rd.w_ptr_r [1] ? _02257_ : _02256_;
  assign _02259_ = \bapg_rd.w_ptr_r [2] ? _02258_ : _02255_;
  assign _02260_ = \bapg_rd.w_ptr_r [3] ? _02259_ : _02252_;
  assign _02261_ = \bapg_rd.w_ptr_r [4] ? _02260_ : _02245_;
  assign _02262_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [1] : \MSYNC_1r1w.synth.nz.mem[160] [1];
  assign _02263_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [1] : \MSYNC_1r1w.synth.nz.mem[162] [1];
  assign _02264_ = \bapg_rd.w_ptr_r [1] ? _02263_ : _02262_;
  assign _02265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [1] : \MSYNC_1r1w.synth.nz.mem[164] [1];
  assign _02266_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [1] : \MSYNC_1r1w.synth.nz.mem[166] [1];
  assign _02267_ = \bapg_rd.w_ptr_r [1] ? _02266_ : _02265_;
  assign _02268_ = \bapg_rd.w_ptr_r [2] ? _02267_ : _02264_;
  assign _02269_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [1] : \MSYNC_1r1w.synth.nz.mem[168] [1];
  assign _02270_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [1] : \MSYNC_1r1w.synth.nz.mem[170] [1];
  assign _02271_ = \bapg_rd.w_ptr_r [1] ? _02270_ : _02269_;
  assign _02272_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [1] : \MSYNC_1r1w.synth.nz.mem[172] [1];
  assign _02273_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [1] : \MSYNC_1r1w.synth.nz.mem[174] [1];
  assign _02274_ = \bapg_rd.w_ptr_r [1] ? _02273_ : _02272_;
  assign _02275_ = \bapg_rd.w_ptr_r [2] ? _02274_ : _02271_;
  assign _02276_ = \bapg_rd.w_ptr_r [3] ? _02275_ : _02268_;
  assign _02277_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [1] : \MSYNC_1r1w.synth.nz.mem[176] [1];
  assign _02278_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [1] : \MSYNC_1r1w.synth.nz.mem[178] [1];
  assign _02279_ = \bapg_rd.w_ptr_r [1] ? _02278_ : _02277_;
  assign _02280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [1] : \MSYNC_1r1w.synth.nz.mem[180] [1];
  assign _02281_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [1] : \MSYNC_1r1w.synth.nz.mem[182] [1];
  assign _02282_ = \bapg_rd.w_ptr_r [1] ? _02281_ : _02280_;
  assign _02283_ = \bapg_rd.w_ptr_r [2] ? _02282_ : _02279_;
  assign _02284_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [1] : \MSYNC_1r1w.synth.nz.mem[184] [1];
  assign _02285_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [1] : \MSYNC_1r1w.synth.nz.mem[186] [1];
  assign _02286_ = \bapg_rd.w_ptr_r [1] ? _02285_ : _02284_;
  assign _02287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [1] : \MSYNC_1r1w.synth.nz.mem[188] [1];
  assign _02288_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [1] : \MSYNC_1r1w.synth.nz.mem[190] [1];
  assign _02289_ = \bapg_rd.w_ptr_r [1] ? _02288_ : _02287_;
  assign _02290_ = \bapg_rd.w_ptr_r [2] ? _02289_ : _02286_;
  assign _02291_ = \bapg_rd.w_ptr_r [3] ? _02290_ : _02283_;
  assign _02292_ = \bapg_rd.w_ptr_r [4] ? _02291_ : _02276_;
  assign _02293_ = \bapg_rd.w_ptr_r [5] ? _02292_ : _02261_;
  assign _02294_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [1] : \MSYNC_1r1w.synth.nz.mem[192] [1];
  assign _02295_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [1] : \MSYNC_1r1w.synth.nz.mem[194] [1];
  assign _02296_ = \bapg_rd.w_ptr_r [1] ? _02295_ : _02294_;
  assign _02297_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [1] : \MSYNC_1r1w.synth.nz.mem[196] [1];
  assign _02298_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [1] : \MSYNC_1r1w.synth.nz.mem[198] [1];
  assign _02299_ = \bapg_rd.w_ptr_r [1] ? _02298_ : _02297_;
  assign _02300_ = \bapg_rd.w_ptr_r [2] ? _02299_ : _02296_;
  assign _02301_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [1] : \MSYNC_1r1w.synth.nz.mem[200] [1];
  assign _02302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [1] : \MSYNC_1r1w.synth.nz.mem[202] [1];
  assign _02303_ = \bapg_rd.w_ptr_r [1] ? _02302_ : _02301_;
  assign _02304_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [1] : \MSYNC_1r1w.synth.nz.mem[204] [1];
  assign _02305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [1] : \MSYNC_1r1w.synth.nz.mem[206] [1];
  assign _02306_ = \bapg_rd.w_ptr_r [1] ? _02305_ : _02304_;
  assign _02307_ = \bapg_rd.w_ptr_r [2] ? _02306_ : _02303_;
  assign _02308_ = \bapg_rd.w_ptr_r [3] ? _02307_ : _02300_;
  assign _02309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [1] : \MSYNC_1r1w.synth.nz.mem[208] [1];
  assign _02310_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [1] : \MSYNC_1r1w.synth.nz.mem[210] [1];
  assign _02311_ = \bapg_rd.w_ptr_r [1] ? _02310_ : _02309_;
  assign _02312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [1] : \MSYNC_1r1w.synth.nz.mem[212] [1];
  assign _02313_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [1] : \MSYNC_1r1w.synth.nz.mem[214] [1];
  assign _02314_ = \bapg_rd.w_ptr_r [1] ? _02313_ : _02312_;
  assign _02315_ = \bapg_rd.w_ptr_r [2] ? _02314_ : _02311_;
  assign _02316_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [1] : \MSYNC_1r1w.synth.nz.mem[216] [1];
  assign _02317_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [1] : \MSYNC_1r1w.synth.nz.mem[218] [1];
  assign _02318_ = \bapg_rd.w_ptr_r [1] ? _02317_ : _02316_;
  assign _02319_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [1] : \MSYNC_1r1w.synth.nz.mem[220] [1];
  assign _02320_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [1] : \MSYNC_1r1w.synth.nz.mem[222] [1];
  assign _02321_ = \bapg_rd.w_ptr_r [1] ? _02320_ : _02319_;
  assign _02322_ = \bapg_rd.w_ptr_r [2] ? _02321_ : _02318_;
  assign _02323_ = \bapg_rd.w_ptr_r [3] ? _02322_ : _02315_;
  assign _02324_ = \bapg_rd.w_ptr_r [4] ? _02323_ : _02308_;
  assign _02325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [1] : \MSYNC_1r1w.synth.nz.mem[224] [1];
  assign _02326_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [1] : \MSYNC_1r1w.synth.nz.mem[226] [1];
  assign _02327_ = \bapg_rd.w_ptr_r [1] ? _02326_ : _02325_;
  assign _02328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [1] : \MSYNC_1r1w.synth.nz.mem[228] [1];
  assign _02329_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [1] : \MSYNC_1r1w.synth.nz.mem[230] [1];
  assign _02330_ = \bapg_rd.w_ptr_r [1] ? _02329_ : _02328_;
  assign _02331_ = \bapg_rd.w_ptr_r [2] ? _02330_ : _02327_;
  assign _02332_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [1] : \MSYNC_1r1w.synth.nz.mem[232] [1];
  assign _02333_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [1] : \MSYNC_1r1w.synth.nz.mem[234] [1];
  assign _02334_ = \bapg_rd.w_ptr_r [1] ? _02333_ : _02332_;
  assign _02335_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [1] : \MSYNC_1r1w.synth.nz.mem[236] [1];
  assign _02336_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [1] : \MSYNC_1r1w.synth.nz.mem[238] [1];
  assign _02337_ = \bapg_rd.w_ptr_r [1] ? _02336_ : _02335_;
  assign _02338_ = \bapg_rd.w_ptr_r [2] ? _02337_ : _02334_;
  assign _02339_ = \bapg_rd.w_ptr_r [3] ? _02338_ : _02331_;
  assign _02340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [1] : \MSYNC_1r1w.synth.nz.mem[240] [1];
  assign _02341_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [1] : \MSYNC_1r1w.synth.nz.mem[242] [1];
  assign _02342_ = \bapg_rd.w_ptr_r [1] ? _02341_ : _02340_;
  assign _02343_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [1] : \MSYNC_1r1w.synth.nz.mem[244] [1];
  assign _02344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [1] : \MSYNC_1r1w.synth.nz.mem[246] [1];
  assign _02345_ = \bapg_rd.w_ptr_r [1] ? _02344_ : _02343_;
  assign _02346_ = \bapg_rd.w_ptr_r [2] ? _02345_ : _02342_;
  assign _02347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [1] : \MSYNC_1r1w.synth.nz.mem[248] [1];
  assign _02348_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [1] : \MSYNC_1r1w.synth.nz.mem[250] [1];
  assign _02349_ = \bapg_rd.w_ptr_r [1] ? _02348_ : _02347_;
  assign _02350_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [1] : \MSYNC_1r1w.synth.nz.mem[252] [1];
  assign _02351_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [1] : \MSYNC_1r1w.synth.nz.mem[254] [1];
  assign _02352_ = \bapg_rd.w_ptr_r [1] ? _02351_ : _02350_;
  assign _02353_ = \bapg_rd.w_ptr_r [2] ? _02352_ : _02349_;
  assign _02354_ = \bapg_rd.w_ptr_r [3] ? _02353_ : _02346_;
  assign _02355_ = \bapg_rd.w_ptr_r [4] ? _02354_ : _02339_;
  assign _02356_ = \bapg_rd.w_ptr_r [5] ? _02355_ : _02324_;
  assign _02357_ = \bapg_rd.w_ptr_r [6] ? _02356_ : _02293_;
  assign _02358_ = \bapg_rd.w_ptr_r [7] ? _02357_ : _02230_;
  assign _02359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [1] : \MSYNC_1r1w.synth.nz.mem[256] [1];
  assign _02360_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [1] : \MSYNC_1r1w.synth.nz.mem[258] [1];
  assign _02361_ = \bapg_rd.w_ptr_r [1] ? _02360_ : _02359_;
  assign _02362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [1] : \MSYNC_1r1w.synth.nz.mem[260] [1];
  assign _02363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [1] : \MSYNC_1r1w.synth.nz.mem[262] [1];
  assign _02364_ = \bapg_rd.w_ptr_r [1] ? _02363_ : _02362_;
  assign _02365_ = \bapg_rd.w_ptr_r [2] ? _02364_ : _02361_;
  assign _02366_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [1] : \MSYNC_1r1w.synth.nz.mem[264] [1];
  assign _02367_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [1] : \MSYNC_1r1w.synth.nz.mem[266] [1];
  assign _02368_ = \bapg_rd.w_ptr_r [1] ? _02367_ : _02366_;
  assign _02369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [1] : \MSYNC_1r1w.synth.nz.mem[268] [1];
  assign _02370_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [1] : \MSYNC_1r1w.synth.nz.mem[270] [1];
  assign _02371_ = \bapg_rd.w_ptr_r [1] ? _02370_ : _02369_;
  assign _02372_ = \bapg_rd.w_ptr_r [2] ? _02371_ : _02368_;
  assign _02373_ = \bapg_rd.w_ptr_r [3] ? _02372_ : _02365_;
  assign _02374_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [1] : \MSYNC_1r1w.synth.nz.mem[272] [1];
  assign _02375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [1] : \MSYNC_1r1w.synth.nz.mem[274] [1];
  assign _02376_ = \bapg_rd.w_ptr_r [1] ? _02375_ : _02374_;
  assign _02377_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [1] : \MSYNC_1r1w.synth.nz.mem[276] [1];
  assign _02378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [1] : \MSYNC_1r1w.synth.nz.mem[278] [1];
  assign _02379_ = \bapg_rd.w_ptr_r [1] ? _02378_ : _02377_;
  assign _02380_ = \bapg_rd.w_ptr_r [2] ? _02379_ : _02376_;
  assign _02381_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [1] : \MSYNC_1r1w.synth.nz.mem[280] [1];
  assign _02382_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [1] : \MSYNC_1r1w.synth.nz.mem[282] [1];
  assign _02383_ = \bapg_rd.w_ptr_r [1] ? _02382_ : _02381_;
  assign _02384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [1] : \MSYNC_1r1w.synth.nz.mem[284] [1];
  assign _02385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [1] : \MSYNC_1r1w.synth.nz.mem[286] [1];
  assign _02386_ = \bapg_rd.w_ptr_r [1] ? _02385_ : _02384_;
  assign _02387_ = \bapg_rd.w_ptr_r [2] ? _02386_ : _02383_;
  assign _02388_ = \bapg_rd.w_ptr_r [3] ? _02387_ : _02380_;
  assign _02389_ = \bapg_rd.w_ptr_r [4] ? _02388_ : _02373_;
  assign _02390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [1] : \MSYNC_1r1w.synth.nz.mem[288] [1];
  assign _02391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [1] : \MSYNC_1r1w.synth.nz.mem[290] [1];
  assign _02392_ = \bapg_rd.w_ptr_r [1] ? _02391_ : _02390_;
  assign _02393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [1] : \MSYNC_1r1w.synth.nz.mem[292] [1];
  assign _02394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [1] : \MSYNC_1r1w.synth.nz.mem[294] [1];
  assign _02395_ = \bapg_rd.w_ptr_r [1] ? _02394_ : _02393_;
  assign _02396_ = \bapg_rd.w_ptr_r [2] ? _02395_ : _02392_;
  assign _02397_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [1] : \MSYNC_1r1w.synth.nz.mem[296] [1];
  assign _02398_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [1] : \MSYNC_1r1w.synth.nz.mem[298] [1];
  assign _02399_ = \bapg_rd.w_ptr_r [1] ? _02398_ : _02397_;
  assign _02400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [1] : \MSYNC_1r1w.synth.nz.mem[300] [1];
  assign _02401_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [1] : \MSYNC_1r1w.synth.nz.mem[302] [1];
  assign _02402_ = \bapg_rd.w_ptr_r [1] ? _02401_ : _02400_;
  assign _02403_ = \bapg_rd.w_ptr_r [2] ? _02402_ : _02399_;
  assign _02404_ = \bapg_rd.w_ptr_r [3] ? _02403_ : _02396_;
  assign _02405_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [1] : \MSYNC_1r1w.synth.nz.mem[304] [1];
  assign _02406_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [1] : \MSYNC_1r1w.synth.nz.mem[306] [1];
  assign _02407_ = \bapg_rd.w_ptr_r [1] ? _02406_ : _02405_;
  assign _02408_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [1] : \MSYNC_1r1w.synth.nz.mem[308] [1];
  assign _02409_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [1] : \MSYNC_1r1w.synth.nz.mem[310] [1];
  assign _02410_ = \bapg_rd.w_ptr_r [1] ? _02409_ : _02408_;
  assign _02411_ = \bapg_rd.w_ptr_r [2] ? _02410_ : _02407_;
  assign _02412_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [1] : \MSYNC_1r1w.synth.nz.mem[312] [1];
  assign _02413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [1] : \MSYNC_1r1w.synth.nz.mem[314] [1];
  assign _02414_ = \bapg_rd.w_ptr_r [1] ? _02413_ : _02412_;
  assign _02415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [1] : \MSYNC_1r1w.synth.nz.mem[316] [1];
  assign _02416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [1] : \MSYNC_1r1w.synth.nz.mem[318] [1];
  assign _02417_ = \bapg_rd.w_ptr_r [1] ? _02416_ : _02415_;
  assign _02418_ = \bapg_rd.w_ptr_r [2] ? _02417_ : _02414_;
  assign _02419_ = \bapg_rd.w_ptr_r [3] ? _02418_ : _02411_;
  assign _02420_ = \bapg_rd.w_ptr_r [4] ? _02419_ : _02404_;
  assign _02421_ = \bapg_rd.w_ptr_r [5] ? _02420_ : _02389_;
  assign _02422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [1] : \MSYNC_1r1w.synth.nz.mem[320] [1];
  assign _02423_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [1] : \MSYNC_1r1w.synth.nz.mem[322] [1];
  assign _02424_ = \bapg_rd.w_ptr_r [1] ? _02423_ : _02422_;
  assign _02425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [1] : \MSYNC_1r1w.synth.nz.mem[324] [1];
  assign _02426_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [1] : \MSYNC_1r1w.synth.nz.mem[326] [1];
  assign _02427_ = \bapg_rd.w_ptr_r [1] ? _02426_ : _02425_;
  assign _02428_ = \bapg_rd.w_ptr_r [2] ? _02427_ : _02424_;
  assign _02429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [1] : \MSYNC_1r1w.synth.nz.mem[328] [1];
  assign _02430_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [1] : \MSYNC_1r1w.synth.nz.mem[330] [1];
  assign _02431_ = \bapg_rd.w_ptr_r [1] ? _02430_ : _02429_;
  assign _02432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [1] : \MSYNC_1r1w.synth.nz.mem[332] [1];
  assign _02433_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [1] : \MSYNC_1r1w.synth.nz.mem[334] [1];
  assign _02434_ = \bapg_rd.w_ptr_r [1] ? _02433_ : _02432_;
  assign _02435_ = \bapg_rd.w_ptr_r [2] ? _02434_ : _02431_;
  assign _02436_ = \bapg_rd.w_ptr_r [3] ? _02435_ : _02428_;
  assign _02437_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [1] : \MSYNC_1r1w.synth.nz.mem[336] [1];
  assign _02438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [1] : \MSYNC_1r1w.synth.nz.mem[338] [1];
  assign _02439_ = \bapg_rd.w_ptr_r [1] ? _02438_ : _02437_;
  assign _02440_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [1] : \MSYNC_1r1w.synth.nz.mem[340] [1];
  assign _02441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [1] : \MSYNC_1r1w.synth.nz.mem[342] [1];
  assign _02442_ = \bapg_rd.w_ptr_r [1] ? _02441_ : _02440_;
  assign _02443_ = \bapg_rd.w_ptr_r [2] ? _02442_ : _02439_;
  assign _02444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [1] : \MSYNC_1r1w.synth.nz.mem[344] [1];
  assign _02445_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [1] : \MSYNC_1r1w.synth.nz.mem[346] [1];
  assign _02446_ = \bapg_rd.w_ptr_r [1] ? _02445_ : _02444_;
  assign _02447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [1] : \MSYNC_1r1w.synth.nz.mem[348] [1];
  assign _02448_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [1] : \MSYNC_1r1w.synth.nz.mem[350] [1];
  assign _02449_ = \bapg_rd.w_ptr_r [1] ? _02448_ : _02447_;
  assign _02450_ = \bapg_rd.w_ptr_r [2] ? _02449_ : _02446_;
  assign _02451_ = \bapg_rd.w_ptr_r [3] ? _02450_ : _02443_;
  assign _02452_ = \bapg_rd.w_ptr_r [4] ? _02451_ : _02436_;
  assign _02453_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [1] : \MSYNC_1r1w.synth.nz.mem[352] [1];
  assign _02454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [1] : \MSYNC_1r1w.synth.nz.mem[354] [1];
  assign _02455_ = \bapg_rd.w_ptr_r [1] ? _02454_ : _02453_;
  assign _02456_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [1] : \MSYNC_1r1w.synth.nz.mem[356] [1];
  assign _02457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [1] : \MSYNC_1r1w.synth.nz.mem[358] [1];
  assign _02458_ = \bapg_rd.w_ptr_r [1] ? _02457_ : _02456_;
  assign _02459_ = \bapg_rd.w_ptr_r [2] ? _02458_ : _02455_;
  assign _02460_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [1] : \MSYNC_1r1w.synth.nz.mem[360] [1];
  assign _02461_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [1] : \MSYNC_1r1w.synth.nz.mem[362] [1];
  assign _02462_ = \bapg_rd.w_ptr_r [1] ? _02461_ : _02460_;
  assign _02463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [1] : \MSYNC_1r1w.synth.nz.mem[364] [1];
  assign _02464_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [1] : \MSYNC_1r1w.synth.nz.mem[366] [1];
  assign _02465_ = \bapg_rd.w_ptr_r [1] ? _02464_ : _02463_;
  assign _02466_ = \bapg_rd.w_ptr_r [2] ? _02465_ : _02462_;
  assign _02467_ = \bapg_rd.w_ptr_r [3] ? _02466_ : _02459_;
  assign _02468_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [1] : \MSYNC_1r1w.synth.nz.mem[368] [1];
  assign _02469_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [1] : \MSYNC_1r1w.synth.nz.mem[370] [1];
  assign _02470_ = \bapg_rd.w_ptr_r [1] ? _02469_ : _02468_;
  assign _02471_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [1] : \MSYNC_1r1w.synth.nz.mem[372] [1];
  assign _02472_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [1] : \MSYNC_1r1w.synth.nz.mem[374] [1];
  assign _02473_ = \bapg_rd.w_ptr_r [1] ? _02472_ : _02471_;
  assign _02474_ = \bapg_rd.w_ptr_r [2] ? _02473_ : _02470_;
  assign _02475_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [1] : \MSYNC_1r1w.synth.nz.mem[376] [1];
  assign _02476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [1] : \MSYNC_1r1w.synth.nz.mem[378] [1];
  assign _02477_ = \bapg_rd.w_ptr_r [1] ? _02476_ : _02475_;
  assign _02478_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [1] : \MSYNC_1r1w.synth.nz.mem[380] [1];
  assign _02479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [1] : \MSYNC_1r1w.synth.nz.mem[382] [1];
  assign _02480_ = \bapg_rd.w_ptr_r [1] ? _02479_ : _02478_;
  assign _02481_ = \bapg_rd.w_ptr_r [2] ? _02480_ : _02477_;
  assign _02482_ = \bapg_rd.w_ptr_r [3] ? _02481_ : _02474_;
  assign _02483_ = \bapg_rd.w_ptr_r [4] ? _02482_ : _02467_;
  assign _02484_ = \bapg_rd.w_ptr_r [5] ? _02483_ : _02452_;
  assign _02485_ = \bapg_rd.w_ptr_r [6] ? _02484_ : _02421_;
  assign _02486_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [1] : \MSYNC_1r1w.synth.nz.mem[384] [1];
  assign _02487_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [1] : \MSYNC_1r1w.synth.nz.mem[386] [1];
  assign _02488_ = \bapg_rd.w_ptr_r [1] ? _02487_ : _02486_;
  assign _02489_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [1] : \MSYNC_1r1w.synth.nz.mem[388] [1];
  assign _02490_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [1] : \MSYNC_1r1w.synth.nz.mem[390] [1];
  assign _02491_ = \bapg_rd.w_ptr_r [1] ? _02490_ : _02489_;
  assign _02492_ = \bapg_rd.w_ptr_r [2] ? _02491_ : _02488_;
  assign _02493_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [1] : \MSYNC_1r1w.synth.nz.mem[392] [1];
  assign _02494_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [1] : \MSYNC_1r1w.synth.nz.mem[394] [1];
  assign _02495_ = \bapg_rd.w_ptr_r [1] ? _02494_ : _02493_;
  assign _02496_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [1] : \MSYNC_1r1w.synth.nz.mem[396] [1];
  assign _02497_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [1] : \MSYNC_1r1w.synth.nz.mem[398] [1];
  assign _02498_ = \bapg_rd.w_ptr_r [1] ? _02497_ : _02496_;
  assign _02499_ = \bapg_rd.w_ptr_r [2] ? _02498_ : _02495_;
  assign _02500_ = \bapg_rd.w_ptr_r [3] ? _02499_ : _02492_;
  assign _02501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [1] : \MSYNC_1r1w.synth.nz.mem[400] [1];
  assign _02502_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [1] : \MSYNC_1r1w.synth.nz.mem[402] [1];
  assign _02503_ = \bapg_rd.w_ptr_r [1] ? _02502_ : _02501_;
  assign _02504_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [1] : \MSYNC_1r1w.synth.nz.mem[404] [1];
  assign _02505_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [1] : \MSYNC_1r1w.synth.nz.mem[406] [1];
  assign _02506_ = \bapg_rd.w_ptr_r [1] ? _02505_ : _02504_;
  assign _02507_ = \bapg_rd.w_ptr_r [2] ? _02506_ : _02503_;
  assign _02508_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [1] : \MSYNC_1r1w.synth.nz.mem[408] [1];
  assign _02509_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [1] : \MSYNC_1r1w.synth.nz.mem[410] [1];
  assign _02510_ = \bapg_rd.w_ptr_r [1] ? _02509_ : _02508_;
  assign _02511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [1] : \MSYNC_1r1w.synth.nz.mem[412] [1];
  assign _02512_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [1] : \MSYNC_1r1w.synth.nz.mem[414] [1];
  assign _02513_ = \bapg_rd.w_ptr_r [1] ? _02512_ : _02511_;
  assign _02514_ = \bapg_rd.w_ptr_r [2] ? _02513_ : _02510_;
  assign _02515_ = \bapg_rd.w_ptr_r [3] ? _02514_ : _02507_;
  assign _02516_ = \bapg_rd.w_ptr_r [4] ? _02515_ : _02500_;
  assign _02517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [1] : \MSYNC_1r1w.synth.nz.mem[416] [1];
  assign _02518_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [1] : \MSYNC_1r1w.synth.nz.mem[418] [1];
  assign _02519_ = \bapg_rd.w_ptr_r [1] ? _02518_ : _02517_;
  assign _02520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [1] : \MSYNC_1r1w.synth.nz.mem[420] [1];
  assign _02521_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [1] : \MSYNC_1r1w.synth.nz.mem[422] [1];
  assign _02522_ = \bapg_rd.w_ptr_r [1] ? _02521_ : _02520_;
  assign _02523_ = \bapg_rd.w_ptr_r [2] ? _02522_ : _02519_;
  assign _02524_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [1] : \MSYNC_1r1w.synth.nz.mem[424] [1];
  assign _02525_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [1] : \MSYNC_1r1w.synth.nz.mem[426] [1];
  assign _02526_ = \bapg_rd.w_ptr_r [1] ? _02525_ : _02524_;
  assign _02527_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [1] : \MSYNC_1r1w.synth.nz.mem[428] [1];
  assign _02528_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [1] : \MSYNC_1r1w.synth.nz.mem[430] [1];
  assign _02529_ = \bapg_rd.w_ptr_r [1] ? _02528_ : _02527_;
  assign _02530_ = \bapg_rd.w_ptr_r [2] ? _02529_ : _02526_;
  assign _02531_ = \bapg_rd.w_ptr_r [3] ? _02530_ : _02523_;
  assign _02532_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [1] : \MSYNC_1r1w.synth.nz.mem[432] [1];
  assign _02533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [1] : \MSYNC_1r1w.synth.nz.mem[434] [1];
  assign _02534_ = \bapg_rd.w_ptr_r [1] ? _02533_ : _02532_;
  assign _02535_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [1] : \MSYNC_1r1w.synth.nz.mem[436] [1];
  assign _02536_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [1] : \MSYNC_1r1w.synth.nz.mem[438] [1];
  assign _02537_ = \bapg_rd.w_ptr_r [1] ? _02536_ : _02535_;
  assign _02538_ = \bapg_rd.w_ptr_r [2] ? _02537_ : _02534_;
  assign _02539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [1] : \MSYNC_1r1w.synth.nz.mem[440] [1];
  assign _02540_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [1] : \MSYNC_1r1w.synth.nz.mem[442] [1];
  assign _02541_ = \bapg_rd.w_ptr_r [1] ? _02540_ : _02539_;
  assign _02542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [1] : \MSYNC_1r1w.synth.nz.mem[444] [1];
  assign _02543_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [1] : \MSYNC_1r1w.synth.nz.mem[446] [1];
  assign _02544_ = \bapg_rd.w_ptr_r [1] ? _02543_ : _02542_;
  assign _02545_ = \bapg_rd.w_ptr_r [2] ? _02544_ : _02541_;
  assign _02546_ = \bapg_rd.w_ptr_r [3] ? _02545_ : _02538_;
  assign _02547_ = \bapg_rd.w_ptr_r [4] ? _02546_ : _02531_;
  assign _02548_ = \bapg_rd.w_ptr_r [5] ? _02547_ : _02516_;
  assign _02549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [1] : \MSYNC_1r1w.synth.nz.mem[448] [1];
  assign _02550_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [1] : \MSYNC_1r1w.synth.nz.mem[450] [1];
  assign _02551_ = \bapg_rd.w_ptr_r [1] ? _02550_ : _02549_;
  assign _02552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [1] : \MSYNC_1r1w.synth.nz.mem[452] [1];
  assign _02553_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [1] : \MSYNC_1r1w.synth.nz.mem[454] [1];
  assign _02554_ = \bapg_rd.w_ptr_r [1] ? _02553_ : _02552_;
  assign _02555_ = \bapg_rd.w_ptr_r [2] ? _02554_ : _02551_;
  assign _02556_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [1] : \MSYNC_1r1w.synth.nz.mem[456] [1];
  assign _02557_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [1] : \MSYNC_1r1w.synth.nz.mem[458] [1];
  assign _02558_ = \bapg_rd.w_ptr_r [1] ? _02557_ : _02556_;
  assign _02559_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [1] : \MSYNC_1r1w.synth.nz.mem[460] [1];
  assign _02560_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [1] : \MSYNC_1r1w.synth.nz.mem[462] [1];
  assign _02561_ = \bapg_rd.w_ptr_r [1] ? _02560_ : _02559_;
  assign _02562_ = \bapg_rd.w_ptr_r [2] ? _02561_ : _02558_;
  assign _02563_ = \bapg_rd.w_ptr_r [3] ? _02562_ : _02555_;
  assign _02564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [1] : \MSYNC_1r1w.synth.nz.mem[464] [1];
  assign _02565_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [1] : \MSYNC_1r1w.synth.nz.mem[466] [1];
  assign _02566_ = \bapg_rd.w_ptr_r [1] ? _02565_ : _02564_;
  assign _02567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [1] : \MSYNC_1r1w.synth.nz.mem[468] [1];
  assign _02568_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [1] : \MSYNC_1r1w.synth.nz.mem[470] [1];
  assign _02569_ = \bapg_rd.w_ptr_r [1] ? _02568_ : _02567_;
  assign _02570_ = \bapg_rd.w_ptr_r [2] ? _02569_ : _02566_;
  assign _02571_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [1] : \MSYNC_1r1w.synth.nz.mem[472] [1];
  assign _02572_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [1] : \MSYNC_1r1w.synth.nz.mem[474] [1];
  assign _02573_ = \bapg_rd.w_ptr_r [1] ? _02572_ : _02571_;
  assign _02574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [1] : \MSYNC_1r1w.synth.nz.mem[476] [1];
  assign _02575_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [1] : \MSYNC_1r1w.synth.nz.mem[478] [1];
  assign _02576_ = \bapg_rd.w_ptr_r [1] ? _02575_ : _02574_;
  assign _02577_ = \bapg_rd.w_ptr_r [2] ? _02576_ : _02573_;
  assign _02578_ = \bapg_rd.w_ptr_r [3] ? _02577_ : _02570_;
  assign _02579_ = \bapg_rd.w_ptr_r [4] ? _02578_ : _02563_;
  assign _02580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [1] : \MSYNC_1r1w.synth.nz.mem[480] [1];
  assign _02581_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [1] : \MSYNC_1r1w.synth.nz.mem[482] [1];
  assign _02582_ = \bapg_rd.w_ptr_r [1] ? _02581_ : _02580_;
  assign _02583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [1] : \MSYNC_1r1w.synth.nz.mem[484] [1];
  assign _02584_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [1] : \MSYNC_1r1w.synth.nz.mem[486] [1];
  assign _02585_ = \bapg_rd.w_ptr_r [1] ? _02584_ : _02583_;
  assign _02586_ = \bapg_rd.w_ptr_r [2] ? _02585_ : _02582_;
  assign _02587_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [1] : \MSYNC_1r1w.synth.nz.mem[488] [1];
  assign _02588_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [1] : \MSYNC_1r1w.synth.nz.mem[490] [1];
  assign _02589_ = \bapg_rd.w_ptr_r [1] ? _02588_ : _02587_;
  assign _02590_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [1] : \MSYNC_1r1w.synth.nz.mem[492] [1];
  assign _02591_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [1] : \MSYNC_1r1w.synth.nz.mem[494] [1];
  assign _02592_ = \bapg_rd.w_ptr_r [1] ? _02591_ : _02590_;
  assign _02593_ = \bapg_rd.w_ptr_r [2] ? _02592_ : _02589_;
  assign _02594_ = \bapg_rd.w_ptr_r [3] ? _02593_ : _02586_;
  assign _02595_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [1] : \MSYNC_1r1w.synth.nz.mem[496] [1];
  assign _02596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [1] : \MSYNC_1r1w.synth.nz.mem[498] [1];
  assign _02597_ = \bapg_rd.w_ptr_r [1] ? _02596_ : _02595_;
  assign _02598_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [1] : \MSYNC_1r1w.synth.nz.mem[500] [1];
  assign _02599_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [1] : \MSYNC_1r1w.synth.nz.mem[502] [1];
  assign _02600_ = \bapg_rd.w_ptr_r [1] ? _02599_ : _02598_;
  assign _02601_ = \bapg_rd.w_ptr_r [2] ? _02600_ : _02597_;
  assign _02602_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [1] : \MSYNC_1r1w.synth.nz.mem[504] [1];
  assign _02603_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [1] : \MSYNC_1r1w.synth.nz.mem[506] [1];
  assign _02604_ = \bapg_rd.w_ptr_r [1] ? _02603_ : _02602_;
  assign _02605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [1] : \MSYNC_1r1w.synth.nz.mem[508] [1];
  assign _02606_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [1] : \MSYNC_1r1w.synth.nz.mem[510] [1];
  assign _02607_ = \bapg_rd.w_ptr_r [1] ? _02606_ : _02605_;
  assign _02608_ = \bapg_rd.w_ptr_r [2] ? _02607_ : _02604_;
  assign _02609_ = \bapg_rd.w_ptr_r [3] ? _02608_ : _02601_;
  assign _02610_ = \bapg_rd.w_ptr_r [4] ? _02609_ : _02594_;
  assign _02611_ = \bapg_rd.w_ptr_r [5] ? _02610_ : _02579_;
  assign _02612_ = \bapg_rd.w_ptr_r [6] ? _02611_ : _02548_;
  assign _02613_ = \bapg_rd.w_ptr_r [7] ? _02612_ : _02485_;
  assign _02614_ = \bapg_rd.w_ptr_r [8] ? _02613_ : _02358_;
  assign _02615_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [1] : \MSYNC_1r1w.synth.nz.mem[512] [1];
  assign _02616_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [1] : \MSYNC_1r1w.synth.nz.mem[514] [1];
  assign _02617_ = \bapg_rd.w_ptr_r [1] ? _02616_ : _02615_;
  assign _02618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [1] : \MSYNC_1r1w.synth.nz.mem[516] [1];
  assign _02619_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [1] : \MSYNC_1r1w.synth.nz.mem[518] [1];
  assign _02620_ = \bapg_rd.w_ptr_r [1] ? _02619_ : _02618_;
  assign _02621_ = \bapg_rd.w_ptr_r [2] ? _02620_ : _02617_;
  assign _02622_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [1] : \MSYNC_1r1w.synth.nz.mem[520] [1];
  assign _02623_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [1] : \MSYNC_1r1w.synth.nz.mem[522] [1];
  assign _02624_ = \bapg_rd.w_ptr_r [1] ? _02623_ : _02622_;
  assign _02625_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [1] : \MSYNC_1r1w.synth.nz.mem[524] [1];
  assign _02626_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [1] : \MSYNC_1r1w.synth.nz.mem[526] [1];
  assign _02627_ = \bapg_rd.w_ptr_r [1] ? _02626_ : _02625_;
  assign _02628_ = \bapg_rd.w_ptr_r [2] ? _02627_ : _02624_;
  assign _02629_ = \bapg_rd.w_ptr_r [3] ? _02628_ : _02621_;
  assign _02630_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [1] : \MSYNC_1r1w.synth.nz.mem[528] [1];
  assign _02631_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [1] : \MSYNC_1r1w.synth.nz.mem[530] [1];
  assign _02632_ = \bapg_rd.w_ptr_r [1] ? _02631_ : _02630_;
  assign _02633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [1] : \MSYNC_1r1w.synth.nz.mem[532] [1];
  assign _02634_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [1] : \MSYNC_1r1w.synth.nz.mem[534] [1];
  assign _02635_ = \bapg_rd.w_ptr_r [1] ? _02634_ : _02633_;
  assign _02636_ = \bapg_rd.w_ptr_r [2] ? _02635_ : _02632_;
  assign _02637_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [1] : \MSYNC_1r1w.synth.nz.mem[536] [1];
  assign _02638_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [1] : \MSYNC_1r1w.synth.nz.mem[538] [1];
  assign _02639_ = \bapg_rd.w_ptr_r [1] ? _02638_ : _02637_;
  assign _02640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [1] : \MSYNC_1r1w.synth.nz.mem[540] [1];
  assign _02641_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [1] : \MSYNC_1r1w.synth.nz.mem[542] [1];
  assign _02642_ = \bapg_rd.w_ptr_r [1] ? _02641_ : _02640_;
  assign _02643_ = \bapg_rd.w_ptr_r [2] ? _02642_ : _02639_;
  assign _02644_ = \bapg_rd.w_ptr_r [3] ? _02643_ : _02636_;
  assign _02645_ = \bapg_rd.w_ptr_r [4] ? _02644_ : _02629_;
  assign _02646_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [1] : \MSYNC_1r1w.synth.nz.mem[544] [1];
  assign _02647_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [1] : \MSYNC_1r1w.synth.nz.mem[546] [1];
  assign _02648_ = \bapg_rd.w_ptr_r [1] ? _02647_ : _02646_;
  assign _02649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [1] : \MSYNC_1r1w.synth.nz.mem[548] [1];
  assign _02650_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [1] : \MSYNC_1r1w.synth.nz.mem[550] [1];
  assign _02651_ = \bapg_rd.w_ptr_r [1] ? _02650_ : _02649_;
  assign _02652_ = \bapg_rd.w_ptr_r [2] ? _02651_ : _02648_;
  assign _02653_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [1] : \MSYNC_1r1w.synth.nz.mem[552] [1];
  assign _02654_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [1] : \MSYNC_1r1w.synth.nz.mem[554] [1];
  assign _02655_ = \bapg_rd.w_ptr_r [1] ? _02654_ : _02653_;
  assign _02656_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [1] : \MSYNC_1r1w.synth.nz.mem[556] [1];
  assign _02657_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [1] : \MSYNC_1r1w.synth.nz.mem[558] [1];
  assign _02658_ = \bapg_rd.w_ptr_r [1] ? _02657_ : _02656_;
  assign _02659_ = \bapg_rd.w_ptr_r [2] ? _02658_ : _02655_;
  assign _02660_ = \bapg_rd.w_ptr_r [3] ? _02659_ : _02652_;
  assign _02661_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [1] : \MSYNC_1r1w.synth.nz.mem[560] [1];
  assign _02662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [1] : \MSYNC_1r1w.synth.nz.mem[562] [1];
  assign _02663_ = \bapg_rd.w_ptr_r [1] ? _02662_ : _02661_;
  assign _02664_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [1] : \MSYNC_1r1w.synth.nz.mem[564] [1];
  assign _02665_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [1] : \MSYNC_1r1w.synth.nz.mem[566] [1];
  assign _02666_ = \bapg_rd.w_ptr_r [1] ? _02665_ : _02664_;
  assign _02667_ = \bapg_rd.w_ptr_r [2] ? _02666_ : _02663_;
  assign _02668_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [1] : \MSYNC_1r1w.synth.nz.mem[568] [1];
  assign _02669_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [1] : \MSYNC_1r1w.synth.nz.mem[570] [1];
  assign _02670_ = \bapg_rd.w_ptr_r [1] ? _02669_ : _02668_;
  assign _02671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [1] : \MSYNC_1r1w.synth.nz.mem[572] [1];
  assign _02672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [1] : \MSYNC_1r1w.synth.nz.mem[574] [1];
  assign _02673_ = \bapg_rd.w_ptr_r [1] ? _02672_ : _02671_;
  assign _02674_ = \bapg_rd.w_ptr_r [2] ? _02673_ : _02670_;
  assign _02675_ = \bapg_rd.w_ptr_r [3] ? _02674_ : _02667_;
  assign _02676_ = \bapg_rd.w_ptr_r [4] ? _02675_ : _02660_;
  assign _02677_ = \bapg_rd.w_ptr_r [5] ? _02676_ : _02645_;
  assign _02678_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [1] : \MSYNC_1r1w.synth.nz.mem[576] [1];
  assign _02679_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [1] : \MSYNC_1r1w.synth.nz.mem[578] [1];
  assign _02680_ = \bapg_rd.w_ptr_r [1] ? _02679_ : _02678_;
  assign _02681_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [1] : \MSYNC_1r1w.synth.nz.mem[580] [1];
  assign _02682_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [1] : \MSYNC_1r1w.synth.nz.mem[582] [1];
  assign _02683_ = \bapg_rd.w_ptr_r [1] ? _02682_ : _02681_;
  assign _02684_ = \bapg_rd.w_ptr_r [2] ? _02683_ : _02680_;
  assign _02685_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [1] : \MSYNC_1r1w.synth.nz.mem[584] [1];
  assign _02686_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [1] : \MSYNC_1r1w.synth.nz.mem[586] [1];
  assign _02687_ = \bapg_rd.w_ptr_r [1] ? _02686_ : _02685_;
  assign _02688_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [1] : \MSYNC_1r1w.synth.nz.mem[588] [1];
  assign _02689_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [1] : \MSYNC_1r1w.synth.nz.mem[590] [1];
  assign _02690_ = \bapg_rd.w_ptr_r [1] ? _02689_ : _02688_;
  assign _02691_ = \bapg_rd.w_ptr_r [2] ? _02690_ : _02687_;
  assign _02692_ = \bapg_rd.w_ptr_r [3] ? _02691_ : _02684_;
  assign _02693_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [1] : \MSYNC_1r1w.synth.nz.mem[592] [1];
  assign _02694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [1] : \MSYNC_1r1w.synth.nz.mem[594] [1];
  assign _02695_ = \bapg_rd.w_ptr_r [1] ? _02694_ : _02693_;
  assign _02696_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [1] : \MSYNC_1r1w.synth.nz.mem[596] [1];
  assign _02697_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [1] : \MSYNC_1r1w.synth.nz.mem[598] [1];
  assign _02698_ = \bapg_rd.w_ptr_r [1] ? _02697_ : _02696_;
  assign _02699_ = \bapg_rd.w_ptr_r [2] ? _02698_ : _02695_;
  assign _02700_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [1] : \MSYNC_1r1w.synth.nz.mem[600] [1];
  assign _02701_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [1] : \MSYNC_1r1w.synth.nz.mem[602] [1];
  assign _02702_ = \bapg_rd.w_ptr_r [1] ? _02701_ : _02700_;
  assign _02703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [1] : \MSYNC_1r1w.synth.nz.mem[604] [1];
  assign _02704_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [1] : \MSYNC_1r1w.synth.nz.mem[606] [1];
  assign _02705_ = \bapg_rd.w_ptr_r [1] ? _02704_ : _02703_;
  assign _02706_ = \bapg_rd.w_ptr_r [2] ? _02705_ : _02702_;
  assign _02707_ = \bapg_rd.w_ptr_r [3] ? _02706_ : _02699_;
  assign _02708_ = \bapg_rd.w_ptr_r [4] ? _02707_ : _02692_;
  assign _02709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [1] : \MSYNC_1r1w.synth.nz.mem[608] [1];
  assign _02710_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [1] : \MSYNC_1r1w.synth.nz.mem[610] [1];
  assign _02711_ = \bapg_rd.w_ptr_r [1] ? _02710_ : _02709_;
  assign _02712_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [1] : \MSYNC_1r1w.synth.nz.mem[612] [1];
  assign _02713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [1] : \MSYNC_1r1w.synth.nz.mem[614] [1];
  assign _02714_ = \bapg_rd.w_ptr_r [1] ? _02713_ : _02712_;
  assign _02715_ = \bapg_rd.w_ptr_r [2] ? _02714_ : _02711_;
  assign _02716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [1] : \MSYNC_1r1w.synth.nz.mem[616] [1];
  assign _02717_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [1] : \MSYNC_1r1w.synth.nz.mem[618] [1];
  assign _02718_ = \bapg_rd.w_ptr_r [1] ? _02717_ : _02716_;
  assign _02719_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [1] : \MSYNC_1r1w.synth.nz.mem[620] [1];
  assign _02720_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [1] : \MSYNC_1r1w.synth.nz.mem[622] [1];
  assign _02721_ = \bapg_rd.w_ptr_r [1] ? _02720_ : _02719_;
  assign _02722_ = \bapg_rd.w_ptr_r [2] ? _02721_ : _02718_;
  assign _02723_ = \bapg_rd.w_ptr_r [3] ? _02722_ : _02715_;
  assign _02724_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [1] : \MSYNC_1r1w.synth.nz.mem[624] [1];
  assign _02725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [1] : \MSYNC_1r1w.synth.nz.mem[626] [1];
  assign _02726_ = \bapg_rd.w_ptr_r [1] ? _02725_ : _02724_;
  assign _02727_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [1] : \MSYNC_1r1w.synth.nz.mem[628] [1];
  assign _02728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [1] : \MSYNC_1r1w.synth.nz.mem[630] [1];
  assign _02729_ = \bapg_rd.w_ptr_r [1] ? _02728_ : _02727_;
  assign _02730_ = \bapg_rd.w_ptr_r [2] ? _02729_ : _02726_;
  assign _02731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [1] : \MSYNC_1r1w.synth.nz.mem[632] [1];
  assign _02732_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [1] : \MSYNC_1r1w.synth.nz.mem[634] [1];
  assign _02733_ = \bapg_rd.w_ptr_r [1] ? _02732_ : _02731_;
  assign _02734_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [1] : \MSYNC_1r1w.synth.nz.mem[636] [1];
  assign _02735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [1] : \MSYNC_1r1w.synth.nz.mem[638] [1];
  assign _02736_ = \bapg_rd.w_ptr_r [1] ? _02735_ : _02734_;
  assign _02737_ = \bapg_rd.w_ptr_r [2] ? _02736_ : _02733_;
  assign _02738_ = \bapg_rd.w_ptr_r [3] ? _02737_ : _02730_;
  assign _02739_ = \bapg_rd.w_ptr_r [4] ? _02738_ : _02723_;
  assign _02740_ = \bapg_rd.w_ptr_r [5] ? _02739_ : _02708_;
  assign _02741_ = \bapg_rd.w_ptr_r [6] ? _02740_ : _02677_;
  assign _02742_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [1] : \MSYNC_1r1w.synth.nz.mem[640] [1];
  assign _02743_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [1] : \MSYNC_1r1w.synth.nz.mem[642] [1];
  assign _02744_ = \bapg_rd.w_ptr_r [1] ? _02743_ : _02742_;
  assign _02745_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [1] : \MSYNC_1r1w.synth.nz.mem[644] [1];
  assign _02746_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [1] : \MSYNC_1r1w.synth.nz.mem[646] [1];
  assign _02747_ = \bapg_rd.w_ptr_r [1] ? _02746_ : _02745_;
  assign _02748_ = \bapg_rd.w_ptr_r [2] ? _02747_ : _02744_;
  assign _02749_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [1] : \MSYNC_1r1w.synth.nz.mem[648] [1];
  assign _02750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [1] : \MSYNC_1r1w.synth.nz.mem[650] [1];
  assign _02751_ = \bapg_rd.w_ptr_r [1] ? _02750_ : _02749_;
  assign _02752_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [1] : \MSYNC_1r1w.synth.nz.mem[652] [1];
  assign _02753_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [1] : \MSYNC_1r1w.synth.nz.mem[654] [1];
  assign _02754_ = \bapg_rd.w_ptr_r [1] ? _02753_ : _02752_;
  assign _02755_ = \bapg_rd.w_ptr_r [2] ? _02754_ : _02751_;
  assign _02756_ = \bapg_rd.w_ptr_r [3] ? _02755_ : _02748_;
  assign _02757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [1] : \MSYNC_1r1w.synth.nz.mem[656] [1];
  assign _02758_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [1] : \MSYNC_1r1w.synth.nz.mem[658] [1];
  assign _02759_ = \bapg_rd.w_ptr_r [1] ? _02758_ : _02757_;
  assign _02760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [1] : \MSYNC_1r1w.synth.nz.mem[660] [1];
  assign _02761_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [1] : \MSYNC_1r1w.synth.nz.mem[662] [1];
  assign _02762_ = \bapg_rd.w_ptr_r [1] ? _02761_ : _02760_;
  assign _02763_ = \bapg_rd.w_ptr_r [2] ? _02762_ : _02759_;
  assign _02764_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [1] : \MSYNC_1r1w.synth.nz.mem[664] [1];
  assign _02765_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [1] : \MSYNC_1r1w.synth.nz.mem[666] [1];
  assign _02766_ = \bapg_rd.w_ptr_r [1] ? _02765_ : _02764_;
  assign _02767_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [1] : \MSYNC_1r1w.synth.nz.mem[668] [1];
  assign _02768_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [1] : \MSYNC_1r1w.synth.nz.mem[670] [1];
  assign _02769_ = \bapg_rd.w_ptr_r [1] ? _02768_ : _02767_;
  assign _02770_ = \bapg_rd.w_ptr_r [2] ? _02769_ : _02766_;
  assign _02771_ = \bapg_rd.w_ptr_r [3] ? _02770_ : _02763_;
  assign _02772_ = \bapg_rd.w_ptr_r [4] ? _02771_ : _02756_;
  assign _02773_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [1] : \MSYNC_1r1w.synth.nz.mem[672] [1];
  assign _02774_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [1] : \MSYNC_1r1w.synth.nz.mem[674] [1];
  assign _02775_ = \bapg_rd.w_ptr_r [1] ? _02774_ : _02773_;
  assign _02776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [1] : \MSYNC_1r1w.synth.nz.mem[676] [1];
  assign _02777_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [1] : \MSYNC_1r1w.synth.nz.mem[678] [1];
  assign _02778_ = \bapg_rd.w_ptr_r [1] ? _02777_ : _02776_;
  assign _02779_ = \bapg_rd.w_ptr_r [2] ? _02778_ : _02775_;
  assign _02780_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [1] : \MSYNC_1r1w.synth.nz.mem[680] [1];
  assign _02781_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [1] : \MSYNC_1r1w.synth.nz.mem[682] [1];
  assign _02782_ = \bapg_rd.w_ptr_r [1] ? _02781_ : _02780_;
  assign _02783_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [1] : \MSYNC_1r1w.synth.nz.mem[684] [1];
  assign _02784_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [1] : \MSYNC_1r1w.synth.nz.mem[686] [1];
  assign _02785_ = \bapg_rd.w_ptr_r [1] ? _02784_ : _02783_;
  assign _02786_ = \bapg_rd.w_ptr_r [2] ? _02785_ : _02782_;
  assign _02787_ = \bapg_rd.w_ptr_r [3] ? _02786_ : _02779_;
  assign _02788_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [1] : \MSYNC_1r1w.synth.nz.mem[688] [1];
  assign _02789_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [1] : \MSYNC_1r1w.synth.nz.mem[690] [1];
  assign _02790_ = \bapg_rd.w_ptr_r [1] ? _02789_ : _02788_;
  assign _02791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [1] : \MSYNC_1r1w.synth.nz.mem[692] [1];
  assign _02792_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [1] : \MSYNC_1r1w.synth.nz.mem[694] [1];
  assign _02793_ = \bapg_rd.w_ptr_r [1] ? _02792_ : _02791_;
  assign _02794_ = \bapg_rd.w_ptr_r [2] ? _02793_ : _02790_;
  assign _02795_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [1] : \MSYNC_1r1w.synth.nz.mem[696] [1];
  assign _02796_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [1] : \MSYNC_1r1w.synth.nz.mem[698] [1];
  assign _02797_ = \bapg_rd.w_ptr_r [1] ? _02796_ : _02795_;
  assign _02798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [1] : \MSYNC_1r1w.synth.nz.mem[700] [1];
  assign _02799_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [1] : \MSYNC_1r1w.synth.nz.mem[702] [1];
  assign _02800_ = \bapg_rd.w_ptr_r [1] ? _02799_ : _02798_;
  assign _02801_ = \bapg_rd.w_ptr_r [2] ? _02800_ : _02797_;
  assign _02802_ = \bapg_rd.w_ptr_r [3] ? _02801_ : _02794_;
  assign _02803_ = \bapg_rd.w_ptr_r [4] ? _02802_ : _02787_;
  assign _02804_ = \bapg_rd.w_ptr_r [5] ? _02803_ : _02772_;
  assign _02805_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [1] : \MSYNC_1r1w.synth.nz.mem[704] [1];
  assign _02806_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [1] : \MSYNC_1r1w.synth.nz.mem[706] [1];
  assign _02807_ = \bapg_rd.w_ptr_r [1] ? _02806_ : _02805_;
  assign _02808_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [1] : \MSYNC_1r1w.synth.nz.mem[708] [1];
  assign _02809_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [1] : \MSYNC_1r1w.synth.nz.mem[710] [1];
  assign _02810_ = \bapg_rd.w_ptr_r [1] ? _02809_ : _02808_;
  assign _02811_ = \bapg_rd.w_ptr_r [2] ? _02810_ : _02807_;
  assign _02812_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [1] : \MSYNC_1r1w.synth.nz.mem[712] [1];
  assign _02813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [1] : \MSYNC_1r1w.synth.nz.mem[714] [1];
  assign _02814_ = \bapg_rd.w_ptr_r [1] ? _02813_ : _02812_;
  assign _02815_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [1] : \MSYNC_1r1w.synth.nz.mem[716] [1];
  assign _02816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [1] : \MSYNC_1r1w.synth.nz.mem[718] [1];
  assign _02817_ = \bapg_rd.w_ptr_r [1] ? _02816_ : _02815_;
  assign _02818_ = \bapg_rd.w_ptr_r [2] ? _02817_ : _02814_;
  assign _02819_ = \bapg_rd.w_ptr_r [3] ? _02818_ : _02811_;
  assign _02820_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [1] : \MSYNC_1r1w.synth.nz.mem[720] [1];
  assign _02821_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [1] : \MSYNC_1r1w.synth.nz.mem[722] [1];
  assign _02822_ = \bapg_rd.w_ptr_r [1] ? _02821_ : _02820_;
  assign _02823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [1] : \MSYNC_1r1w.synth.nz.mem[724] [1];
  assign _02824_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [1] : \MSYNC_1r1w.synth.nz.mem[726] [1];
  assign _02825_ = \bapg_rd.w_ptr_r [1] ? _02824_ : _02823_;
  assign _02826_ = \bapg_rd.w_ptr_r [2] ? _02825_ : _02822_;
  assign _02827_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [1] : \MSYNC_1r1w.synth.nz.mem[728] [1];
  assign _02828_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [1] : \MSYNC_1r1w.synth.nz.mem[730] [1];
  assign _02829_ = \bapg_rd.w_ptr_r [1] ? _02828_ : _02827_;
  assign _02830_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [1] : \MSYNC_1r1w.synth.nz.mem[732] [1];
  assign _02831_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [1] : \MSYNC_1r1w.synth.nz.mem[734] [1];
  assign _02832_ = \bapg_rd.w_ptr_r [1] ? _02831_ : _02830_;
  assign _02833_ = \bapg_rd.w_ptr_r [2] ? _02832_ : _02829_;
  assign _02834_ = \bapg_rd.w_ptr_r [3] ? _02833_ : _02826_;
  assign _02835_ = \bapg_rd.w_ptr_r [4] ? _02834_ : _02819_;
  assign _02836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [1] : \MSYNC_1r1w.synth.nz.mem[736] [1];
  assign _02837_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [1] : \MSYNC_1r1w.synth.nz.mem[738] [1];
  assign _02838_ = \bapg_rd.w_ptr_r [1] ? _02837_ : _02836_;
  assign _02839_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [1] : \MSYNC_1r1w.synth.nz.mem[740] [1];
  assign _02840_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [1] : \MSYNC_1r1w.synth.nz.mem[742] [1];
  assign _02841_ = \bapg_rd.w_ptr_r [1] ? _02840_ : _02839_;
  assign _02842_ = \bapg_rd.w_ptr_r [2] ? _02841_ : _02838_;
  assign _02843_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [1] : \MSYNC_1r1w.synth.nz.mem[744] [1];
  assign _02844_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [1] : \MSYNC_1r1w.synth.nz.mem[746] [1];
  assign _02845_ = \bapg_rd.w_ptr_r [1] ? _02844_ : _02843_;
  assign _02846_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [1] : \MSYNC_1r1w.synth.nz.mem[748] [1];
  assign _02847_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [1] : \MSYNC_1r1w.synth.nz.mem[750] [1];
  assign _02848_ = \bapg_rd.w_ptr_r [1] ? _02847_ : _02846_;
  assign _02849_ = \bapg_rd.w_ptr_r [2] ? _02848_ : _02845_;
  assign _02850_ = \bapg_rd.w_ptr_r [3] ? _02849_ : _02842_;
  assign _02851_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [1] : \MSYNC_1r1w.synth.nz.mem[752] [1];
  assign _02852_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [1] : \MSYNC_1r1w.synth.nz.mem[754] [1];
  assign _02853_ = \bapg_rd.w_ptr_r [1] ? _02852_ : _02851_;
  assign _02854_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [1] : \MSYNC_1r1w.synth.nz.mem[756] [1];
  assign _02855_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [1] : \MSYNC_1r1w.synth.nz.mem[758] [1];
  assign _02856_ = \bapg_rd.w_ptr_r [1] ? _02855_ : _02854_;
  assign _02857_ = \bapg_rd.w_ptr_r [2] ? _02856_ : _02853_;
  assign _02858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [1] : \MSYNC_1r1w.synth.nz.mem[760] [1];
  assign _02859_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [1] : \MSYNC_1r1w.synth.nz.mem[762] [1];
  assign _02860_ = \bapg_rd.w_ptr_r [1] ? _02859_ : _02858_;
  assign _02861_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [1] : \MSYNC_1r1w.synth.nz.mem[764] [1];
  assign _02862_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [1] : \MSYNC_1r1w.synth.nz.mem[766] [1];
  assign _02863_ = \bapg_rd.w_ptr_r [1] ? _02862_ : _02861_;
  assign _02864_ = \bapg_rd.w_ptr_r [2] ? _02863_ : _02860_;
  assign _02865_ = \bapg_rd.w_ptr_r [3] ? _02864_ : _02857_;
  assign _02866_ = \bapg_rd.w_ptr_r [4] ? _02865_ : _02850_;
  assign _02867_ = \bapg_rd.w_ptr_r [5] ? _02866_ : _02835_;
  assign _02868_ = \bapg_rd.w_ptr_r [6] ? _02867_ : _02804_;
  assign _02869_ = \bapg_rd.w_ptr_r [7] ? _02868_ : _02741_;
  assign _02870_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [1] : \MSYNC_1r1w.synth.nz.mem[768] [1];
  assign _02871_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [1] : \MSYNC_1r1w.synth.nz.mem[770] [1];
  assign _02872_ = \bapg_rd.w_ptr_r [1] ? _02871_ : _02870_;
  assign _02873_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [1] : \MSYNC_1r1w.synth.nz.mem[772] [1];
  assign _02874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [1] : \MSYNC_1r1w.synth.nz.mem[774] [1];
  assign _02875_ = \bapg_rd.w_ptr_r [1] ? _02874_ : _02873_;
  assign _02876_ = \bapg_rd.w_ptr_r [2] ? _02875_ : _02872_;
  assign _02877_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [1] : \MSYNC_1r1w.synth.nz.mem[776] [1];
  assign _02878_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [1] : \MSYNC_1r1w.synth.nz.mem[778] [1];
  assign _02879_ = \bapg_rd.w_ptr_r [1] ? _02878_ : _02877_;
  assign _02880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [1] : \MSYNC_1r1w.synth.nz.mem[780] [1];
  assign _02881_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [1] : \MSYNC_1r1w.synth.nz.mem[782] [1];
  assign _02882_ = \bapg_rd.w_ptr_r [1] ? _02881_ : _02880_;
  assign _02883_ = \bapg_rd.w_ptr_r [2] ? _02882_ : _02879_;
  assign _02884_ = \bapg_rd.w_ptr_r [3] ? _02883_ : _02876_;
  assign _02885_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [1] : \MSYNC_1r1w.synth.nz.mem[784] [1];
  assign _02886_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [1] : \MSYNC_1r1w.synth.nz.mem[786] [1];
  assign _02887_ = \bapg_rd.w_ptr_r [1] ? _02886_ : _02885_;
  assign _02888_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [1] : \MSYNC_1r1w.synth.nz.mem[788] [1];
  assign _02889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [1] : \MSYNC_1r1w.synth.nz.mem[790] [1];
  assign _02890_ = \bapg_rd.w_ptr_r [1] ? _02889_ : _02888_;
  assign _02891_ = \bapg_rd.w_ptr_r [2] ? _02890_ : _02887_;
  assign _02892_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [1] : \MSYNC_1r1w.synth.nz.mem[792] [1];
  assign _02893_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [1] : \MSYNC_1r1w.synth.nz.mem[794] [1];
  assign _02894_ = \bapg_rd.w_ptr_r [1] ? _02893_ : _02892_;
  assign _02895_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [1] : \MSYNC_1r1w.synth.nz.mem[796] [1];
  assign _02896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [1] : \MSYNC_1r1w.synth.nz.mem[798] [1];
  assign _02897_ = \bapg_rd.w_ptr_r [1] ? _02896_ : _02895_;
  assign _02898_ = \bapg_rd.w_ptr_r [2] ? _02897_ : _02894_;
  assign _02899_ = \bapg_rd.w_ptr_r [3] ? _02898_ : _02891_;
  assign _02900_ = \bapg_rd.w_ptr_r [4] ? _02899_ : _02884_;
  assign _02901_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [1] : \MSYNC_1r1w.synth.nz.mem[800] [1];
  assign _02902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [1] : \MSYNC_1r1w.synth.nz.mem[802] [1];
  assign _02903_ = \bapg_rd.w_ptr_r [1] ? _02902_ : _02901_;
  assign _02904_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [1] : \MSYNC_1r1w.synth.nz.mem[804] [1];
  assign _02905_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [1] : \MSYNC_1r1w.synth.nz.mem[806] [1];
  assign _02906_ = \bapg_rd.w_ptr_r [1] ? _02905_ : _02904_;
  assign _02907_ = \bapg_rd.w_ptr_r [2] ? _02906_ : _02903_;
  assign _02908_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [1] : \MSYNC_1r1w.synth.nz.mem[808] [1];
  assign _02909_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [1] : \MSYNC_1r1w.synth.nz.mem[810] [1];
  assign _02910_ = \bapg_rd.w_ptr_r [1] ? _02909_ : _02908_;
  assign _02911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [1] : \MSYNC_1r1w.synth.nz.mem[812] [1];
  assign _02912_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [1] : \MSYNC_1r1w.synth.nz.mem[814] [1];
  assign _02913_ = \bapg_rd.w_ptr_r [1] ? _02912_ : _02911_;
  assign _02914_ = \bapg_rd.w_ptr_r [2] ? _02913_ : _02910_;
  assign _02915_ = \bapg_rd.w_ptr_r [3] ? _02914_ : _02907_;
  assign _02916_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [1] : \MSYNC_1r1w.synth.nz.mem[816] [1];
  assign _02917_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [1] : \MSYNC_1r1w.synth.nz.mem[818] [1];
  assign _02918_ = \bapg_rd.w_ptr_r [1] ? _02917_ : _02916_;
  assign _02919_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [1] : \MSYNC_1r1w.synth.nz.mem[820] [1];
  assign _02920_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [1] : \MSYNC_1r1w.synth.nz.mem[822] [1];
  assign _02921_ = \bapg_rd.w_ptr_r [1] ? _02920_ : _02919_;
  assign _02922_ = \bapg_rd.w_ptr_r [2] ? _02921_ : _02918_;
  assign _02923_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [1] : \MSYNC_1r1w.synth.nz.mem[824] [1];
  assign _02924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [1] : \MSYNC_1r1w.synth.nz.mem[826] [1];
  assign _02925_ = \bapg_rd.w_ptr_r [1] ? _02924_ : _02923_;
  assign _02926_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [1] : \MSYNC_1r1w.synth.nz.mem[828] [1];
  assign _02927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [1] : \MSYNC_1r1w.synth.nz.mem[830] [1];
  assign _02928_ = \bapg_rd.w_ptr_r [1] ? _02927_ : _02926_;
  assign _02929_ = \bapg_rd.w_ptr_r [2] ? _02928_ : _02925_;
  assign _02930_ = \bapg_rd.w_ptr_r [3] ? _02929_ : _02922_;
  assign _02931_ = \bapg_rd.w_ptr_r [4] ? _02930_ : _02915_;
  assign _02932_ = \bapg_rd.w_ptr_r [5] ? _02931_ : _02900_;
  assign _02933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [1] : \MSYNC_1r1w.synth.nz.mem[832] [1];
  assign _02934_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [1] : \MSYNC_1r1w.synth.nz.mem[834] [1];
  assign _02935_ = \bapg_rd.w_ptr_r [1] ? _02934_ : _02933_;
  assign _02936_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [1] : \MSYNC_1r1w.synth.nz.mem[836] [1];
  assign _02937_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [1] : \MSYNC_1r1w.synth.nz.mem[838] [1];
  assign _02938_ = \bapg_rd.w_ptr_r [1] ? _02937_ : _02936_;
  assign _02939_ = \bapg_rd.w_ptr_r [2] ? _02938_ : _02935_;
  assign _02940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [1] : \MSYNC_1r1w.synth.nz.mem[840] [1];
  assign _02941_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [1] : \MSYNC_1r1w.synth.nz.mem[842] [1];
  assign _02942_ = \bapg_rd.w_ptr_r [1] ? _02941_ : _02940_;
  assign _02943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [1] : \MSYNC_1r1w.synth.nz.mem[844] [1];
  assign _02944_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [1] : \MSYNC_1r1w.synth.nz.mem[846] [1];
  assign _02945_ = \bapg_rd.w_ptr_r [1] ? _02944_ : _02943_;
  assign _02946_ = \bapg_rd.w_ptr_r [2] ? _02945_ : _02942_;
  assign _02947_ = \bapg_rd.w_ptr_r [3] ? _02946_ : _02939_;
  assign _02948_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [1] : \MSYNC_1r1w.synth.nz.mem[848] [1];
  assign _02949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [1] : \MSYNC_1r1w.synth.nz.mem[850] [1];
  assign _02950_ = \bapg_rd.w_ptr_r [1] ? _02949_ : _02948_;
  assign _02951_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [1] : \MSYNC_1r1w.synth.nz.mem[852] [1];
  assign _02952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [1] : \MSYNC_1r1w.synth.nz.mem[854] [1];
  assign _02953_ = \bapg_rd.w_ptr_r [1] ? _02952_ : _02951_;
  assign _02954_ = \bapg_rd.w_ptr_r [2] ? _02953_ : _02950_;
  assign _02955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [1] : \MSYNC_1r1w.synth.nz.mem[856] [1];
  assign _02956_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [1] : \MSYNC_1r1w.synth.nz.mem[858] [1];
  assign _02957_ = \bapg_rd.w_ptr_r [1] ? _02956_ : _02955_;
  assign _02958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [1] : \MSYNC_1r1w.synth.nz.mem[860] [1];
  assign _02959_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [1] : \MSYNC_1r1w.synth.nz.mem[862] [1];
  assign _02960_ = \bapg_rd.w_ptr_r [1] ? _02959_ : _02958_;
  assign _02961_ = \bapg_rd.w_ptr_r [2] ? _02960_ : _02957_;
  assign _02962_ = \bapg_rd.w_ptr_r [3] ? _02961_ : _02954_;
  assign _02963_ = \bapg_rd.w_ptr_r [4] ? _02962_ : _02947_;
  assign _02964_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [1] : \MSYNC_1r1w.synth.nz.mem[864] [1];
  assign _02965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [1] : \MSYNC_1r1w.synth.nz.mem[866] [1];
  assign _02966_ = \bapg_rd.w_ptr_r [1] ? _02965_ : _02964_;
  assign _02967_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [1] : \MSYNC_1r1w.synth.nz.mem[868] [1];
  assign _02968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [1] : \MSYNC_1r1w.synth.nz.mem[870] [1];
  assign _02969_ = \bapg_rd.w_ptr_r [1] ? _02968_ : _02967_;
  assign _02970_ = \bapg_rd.w_ptr_r [2] ? _02969_ : _02966_;
  assign _02971_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [1] : \MSYNC_1r1w.synth.nz.mem[872] [1];
  assign _02972_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [1] : \MSYNC_1r1w.synth.nz.mem[874] [1];
  assign _02973_ = \bapg_rd.w_ptr_r [1] ? _02972_ : _02971_;
  assign _02974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [1] : \MSYNC_1r1w.synth.nz.mem[876] [1];
  assign _02975_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [1] : \MSYNC_1r1w.synth.nz.mem[878] [1];
  assign _02976_ = \bapg_rd.w_ptr_r [1] ? _02975_ : _02974_;
  assign _02977_ = \bapg_rd.w_ptr_r [2] ? _02976_ : _02973_;
  assign _02978_ = \bapg_rd.w_ptr_r [3] ? _02977_ : _02970_;
  assign _02979_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [1] : \MSYNC_1r1w.synth.nz.mem[880] [1];
  assign _02980_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [1] : \MSYNC_1r1w.synth.nz.mem[882] [1];
  assign _02981_ = \bapg_rd.w_ptr_r [1] ? _02980_ : _02979_;
  assign _02982_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [1] : \MSYNC_1r1w.synth.nz.mem[884] [1];
  assign _02983_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [1] : \MSYNC_1r1w.synth.nz.mem[886] [1];
  assign _02984_ = \bapg_rd.w_ptr_r [1] ? _02983_ : _02982_;
  assign _02985_ = \bapg_rd.w_ptr_r [2] ? _02984_ : _02981_;
  assign _02986_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [1] : \MSYNC_1r1w.synth.nz.mem[888] [1];
  assign _02987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [1] : \MSYNC_1r1w.synth.nz.mem[890] [1];
  assign _02988_ = \bapg_rd.w_ptr_r [1] ? _02987_ : _02986_;
  assign _02989_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [1] : \MSYNC_1r1w.synth.nz.mem[892] [1];
  assign _02990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [1] : \MSYNC_1r1w.synth.nz.mem[894] [1];
  assign _02991_ = \bapg_rd.w_ptr_r [1] ? _02990_ : _02989_;
  assign _02992_ = \bapg_rd.w_ptr_r [2] ? _02991_ : _02988_;
  assign _02993_ = \bapg_rd.w_ptr_r [3] ? _02992_ : _02985_;
  assign _02994_ = \bapg_rd.w_ptr_r [4] ? _02993_ : _02978_;
  assign _02995_ = \bapg_rd.w_ptr_r [5] ? _02994_ : _02963_;
  assign _02996_ = \bapg_rd.w_ptr_r [6] ? _02995_ : _02932_;
  assign _02997_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [1] : \MSYNC_1r1w.synth.nz.mem[896] [1];
  assign _02998_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [1] : \MSYNC_1r1w.synth.nz.mem[898] [1];
  assign _02999_ = \bapg_rd.w_ptr_r [1] ? _02998_ : _02997_;
  assign _03000_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [1] : \MSYNC_1r1w.synth.nz.mem[900] [1];
  assign _03001_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [1] : \MSYNC_1r1w.synth.nz.mem[902] [1];
  assign _03002_ = \bapg_rd.w_ptr_r [1] ? _03001_ : _03000_;
  assign _03003_ = \bapg_rd.w_ptr_r [2] ? _03002_ : _02999_;
  assign _03004_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [1] : \MSYNC_1r1w.synth.nz.mem[904] [1];
  assign _03005_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [1] : \MSYNC_1r1w.synth.nz.mem[906] [1];
  assign _03006_ = \bapg_rd.w_ptr_r [1] ? _03005_ : _03004_;
  assign _03007_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [1] : \MSYNC_1r1w.synth.nz.mem[908] [1];
  assign _03008_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [1] : \MSYNC_1r1w.synth.nz.mem[910] [1];
  assign _03009_ = \bapg_rd.w_ptr_r [1] ? _03008_ : _03007_;
  assign _03010_ = \bapg_rd.w_ptr_r [2] ? _03009_ : _03006_;
  assign _03011_ = \bapg_rd.w_ptr_r [3] ? _03010_ : _03003_;
  assign _03012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [1] : \MSYNC_1r1w.synth.nz.mem[912] [1];
  assign _03013_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [1] : \MSYNC_1r1w.synth.nz.mem[914] [1];
  assign _03014_ = \bapg_rd.w_ptr_r [1] ? _03013_ : _03012_;
  assign _03015_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [1] : \MSYNC_1r1w.synth.nz.mem[916] [1];
  assign _03016_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [1] : \MSYNC_1r1w.synth.nz.mem[918] [1];
  assign _03017_ = \bapg_rd.w_ptr_r [1] ? _03016_ : _03015_;
  assign _03018_ = \bapg_rd.w_ptr_r [2] ? _03017_ : _03014_;
  assign _03019_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [1] : \MSYNC_1r1w.synth.nz.mem[920] [1];
  assign _03020_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [1] : \MSYNC_1r1w.synth.nz.mem[922] [1];
  assign _03021_ = \bapg_rd.w_ptr_r [1] ? _03020_ : _03019_;
  assign _03022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [1] : \MSYNC_1r1w.synth.nz.mem[924] [1];
  assign _03023_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [1] : \MSYNC_1r1w.synth.nz.mem[926] [1];
  assign _03024_ = \bapg_rd.w_ptr_r [1] ? _03023_ : _03022_;
  assign _03025_ = \bapg_rd.w_ptr_r [2] ? _03024_ : _03021_;
  assign _03026_ = \bapg_rd.w_ptr_r [3] ? _03025_ : _03018_;
  assign _03027_ = \bapg_rd.w_ptr_r [4] ? _03026_ : _03011_;
  assign _03028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [1] : \MSYNC_1r1w.synth.nz.mem[928] [1];
  assign _03029_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [1] : \MSYNC_1r1w.synth.nz.mem[930] [1];
  assign _03030_ = \bapg_rd.w_ptr_r [1] ? _03029_ : _03028_;
  assign _03031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [1] : \MSYNC_1r1w.synth.nz.mem[932] [1];
  assign _03032_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [1] : \MSYNC_1r1w.synth.nz.mem[934] [1];
  assign _03033_ = \bapg_rd.w_ptr_r [1] ? _03032_ : _03031_;
  assign _03034_ = \bapg_rd.w_ptr_r [2] ? _03033_ : _03030_;
  assign _03035_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [1] : \MSYNC_1r1w.synth.nz.mem[936] [1];
  assign _03036_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [1] : \MSYNC_1r1w.synth.nz.mem[938] [1];
  assign _03037_ = \bapg_rd.w_ptr_r [1] ? _03036_ : _03035_;
  assign _03038_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [1] : \MSYNC_1r1w.synth.nz.mem[940] [1];
  assign _03039_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [1] : \MSYNC_1r1w.synth.nz.mem[942] [1];
  assign _03040_ = \bapg_rd.w_ptr_r [1] ? _03039_ : _03038_;
  assign _03041_ = \bapg_rd.w_ptr_r [2] ? _03040_ : _03037_;
  assign _03042_ = \bapg_rd.w_ptr_r [3] ? _03041_ : _03034_;
  assign _03043_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [1] : \MSYNC_1r1w.synth.nz.mem[944] [1];
  assign _03044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [1] : \MSYNC_1r1w.synth.nz.mem[946] [1];
  assign _03045_ = \bapg_rd.w_ptr_r [1] ? _03044_ : _03043_;
  assign _03046_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [1] : \MSYNC_1r1w.synth.nz.mem[948] [1];
  assign _03047_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [1] : \MSYNC_1r1w.synth.nz.mem[950] [1];
  assign _03048_ = \bapg_rd.w_ptr_r [1] ? _03047_ : _03046_;
  assign _03049_ = \bapg_rd.w_ptr_r [2] ? _03048_ : _03045_;
  assign _03050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [1] : \MSYNC_1r1w.synth.nz.mem[952] [1];
  assign _03051_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [1] : \MSYNC_1r1w.synth.nz.mem[954] [1];
  assign _03052_ = \bapg_rd.w_ptr_r [1] ? _03051_ : _03050_;
  assign _03053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [1] : \MSYNC_1r1w.synth.nz.mem[956] [1];
  assign _03054_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [1] : \MSYNC_1r1w.synth.nz.mem[958] [1];
  assign _03055_ = \bapg_rd.w_ptr_r [1] ? _03054_ : _03053_;
  assign _03056_ = \bapg_rd.w_ptr_r [2] ? _03055_ : _03052_;
  assign _03057_ = \bapg_rd.w_ptr_r [3] ? _03056_ : _03049_;
  assign _03058_ = \bapg_rd.w_ptr_r [4] ? _03057_ : _03042_;
  assign _03059_ = \bapg_rd.w_ptr_r [5] ? _03058_ : _03027_;
  assign _03060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [1] : \MSYNC_1r1w.synth.nz.mem[960] [1];
  assign _03061_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [1] : \MSYNC_1r1w.synth.nz.mem[962] [1];
  assign _03062_ = \bapg_rd.w_ptr_r [1] ? _03061_ : _03060_;
  assign _03063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [1] : \MSYNC_1r1w.synth.nz.mem[964] [1];
  assign _03064_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [1] : \MSYNC_1r1w.synth.nz.mem[966] [1];
  assign _03065_ = \bapg_rd.w_ptr_r [1] ? _03064_ : _03063_;
  assign _03066_ = \bapg_rd.w_ptr_r [2] ? _03065_ : _03062_;
  assign _03067_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [1] : \MSYNC_1r1w.synth.nz.mem[968] [1];
  assign _03068_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [1] : \MSYNC_1r1w.synth.nz.mem[970] [1];
  assign _03069_ = \bapg_rd.w_ptr_r [1] ? _03068_ : _03067_;
  assign _03070_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [1] : \MSYNC_1r1w.synth.nz.mem[972] [1];
  assign _03071_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [1] : \MSYNC_1r1w.synth.nz.mem[974] [1];
  assign _03072_ = \bapg_rd.w_ptr_r [1] ? _03071_ : _03070_;
  assign _03073_ = \bapg_rd.w_ptr_r [2] ? _03072_ : _03069_;
  assign _03074_ = \bapg_rd.w_ptr_r [3] ? _03073_ : _03066_;
  assign _03075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [1] : \MSYNC_1r1w.synth.nz.mem[976] [1];
  assign _03076_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [1] : \MSYNC_1r1w.synth.nz.mem[978] [1];
  assign _03077_ = \bapg_rd.w_ptr_r [1] ? _03076_ : _03075_;
  assign _03078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [1] : \MSYNC_1r1w.synth.nz.mem[980] [1];
  assign _03079_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [1] : \MSYNC_1r1w.synth.nz.mem[982] [1];
  assign _03080_ = \bapg_rd.w_ptr_r [1] ? _03079_ : _03078_;
  assign _03081_ = \bapg_rd.w_ptr_r [2] ? _03080_ : _03077_;
  assign _03082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [1] : \MSYNC_1r1w.synth.nz.mem[984] [1];
  assign _03083_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [1] : \MSYNC_1r1w.synth.nz.mem[986] [1];
  assign _03084_ = \bapg_rd.w_ptr_r [1] ? _03083_ : _03082_;
  assign _03085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [1] : \MSYNC_1r1w.synth.nz.mem[988] [1];
  assign _03086_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [1] : \MSYNC_1r1w.synth.nz.mem[990] [1];
  assign _03087_ = \bapg_rd.w_ptr_r [1] ? _03086_ : _03085_;
  assign _03088_ = \bapg_rd.w_ptr_r [2] ? _03087_ : _03084_;
  assign _03089_ = \bapg_rd.w_ptr_r [3] ? _03088_ : _03081_;
  assign _03090_ = \bapg_rd.w_ptr_r [4] ? _03089_ : _03074_;
  assign _03091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [1] : \MSYNC_1r1w.synth.nz.mem[992] [1];
  assign _03092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [1] : \MSYNC_1r1w.synth.nz.mem[994] [1];
  assign _03093_ = \bapg_rd.w_ptr_r [1] ? _03092_ : _03091_;
  assign _03094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [1] : \MSYNC_1r1w.synth.nz.mem[996] [1];
  assign _03095_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [1] : \MSYNC_1r1w.synth.nz.mem[998] [1];
  assign _03096_ = \bapg_rd.w_ptr_r [1] ? _03095_ : _03094_;
  assign _03097_ = \bapg_rd.w_ptr_r [2] ? _03096_ : _03093_;
  assign _03098_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [1] : \MSYNC_1r1w.synth.nz.mem[1000] [1];
  assign _03099_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [1] : \MSYNC_1r1w.synth.nz.mem[1002] [1];
  assign _03100_ = \bapg_rd.w_ptr_r [1] ? _03099_ : _03098_;
  assign _03101_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [1] : \MSYNC_1r1w.synth.nz.mem[1004] [1];
  assign _03102_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [1] : \MSYNC_1r1w.synth.nz.mem[1006] [1];
  assign _03103_ = \bapg_rd.w_ptr_r [1] ? _03102_ : _03101_;
  assign _03104_ = \bapg_rd.w_ptr_r [2] ? _03103_ : _03100_;
  assign _03105_ = \bapg_rd.w_ptr_r [3] ? _03104_ : _03097_;
  assign _03106_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [1] : \MSYNC_1r1w.synth.nz.mem[1008] [1];
  assign _03107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [1] : \MSYNC_1r1w.synth.nz.mem[1010] [1];
  assign _03108_ = \bapg_rd.w_ptr_r [1] ? _03107_ : _03106_;
  assign _03109_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [1] : \MSYNC_1r1w.synth.nz.mem[1012] [1];
  assign _03110_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [1] : \MSYNC_1r1w.synth.nz.mem[1014] [1];
  assign _03111_ = \bapg_rd.w_ptr_r [1] ? _03110_ : _03109_;
  assign _03112_ = \bapg_rd.w_ptr_r [2] ? _03111_ : _03108_;
  assign _03113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [1] : \MSYNC_1r1w.synth.nz.mem[1016] [1];
  assign _03114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [1] : \MSYNC_1r1w.synth.nz.mem[1018] [1];
  assign _03115_ = \bapg_rd.w_ptr_r [1] ? _03114_ : _03113_;
  assign _03116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [1] : \MSYNC_1r1w.synth.nz.mem[1020] [1];
  assign _03117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [1] : \MSYNC_1r1w.synth.nz.mem[1022] [1];
  assign _03118_ = \bapg_rd.w_ptr_r [1] ? _03117_ : _03116_;
  assign _03119_ = \bapg_rd.w_ptr_r [2] ? _03118_ : _03115_;
  assign _03120_ = \bapg_rd.w_ptr_r [3] ? _03119_ : _03112_;
  assign _03121_ = \bapg_rd.w_ptr_r [4] ? _03120_ : _03105_;
  assign _03122_ = \bapg_rd.w_ptr_r [5] ? _03121_ : _03090_;
  assign _03123_ = \bapg_rd.w_ptr_r [6] ? _03122_ : _03059_;
  assign _03124_ = \bapg_rd.w_ptr_r [7] ? _03123_ : _02996_;
  assign _03125_ = \bapg_rd.w_ptr_r [8] ? _03124_ : _02869_;
  assign r_data_o[1] = \bapg_rd.w_ptr_r [9] ? _03125_ : _02614_;
  assign _03126_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [2] : \MSYNC_1r1w.synth.nz.mem[0] [2];
  assign _03127_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [2] : \MSYNC_1r1w.synth.nz.mem[2] [2];
  assign _03128_ = \bapg_rd.w_ptr_r [1] ? _03127_ : _03126_;
  assign _03129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [2] : \MSYNC_1r1w.synth.nz.mem[4] [2];
  assign _03130_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [2] : \MSYNC_1r1w.synth.nz.mem[6] [2];
  assign _03131_ = \bapg_rd.w_ptr_r [1] ? _03130_ : _03129_;
  assign _03132_ = \bapg_rd.w_ptr_r [2] ? _03131_ : _03128_;
  assign _03133_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [2] : \MSYNC_1r1w.synth.nz.mem[8] [2];
  assign _03134_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [2] : \MSYNC_1r1w.synth.nz.mem[10] [2];
  assign _03135_ = \bapg_rd.w_ptr_r [1] ? _03134_ : _03133_;
  assign _03136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [2] : \MSYNC_1r1w.synth.nz.mem[12] [2];
  assign _03137_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [2] : \MSYNC_1r1w.synth.nz.mem[14] [2];
  assign _03138_ = \bapg_rd.w_ptr_r [1] ? _03137_ : _03136_;
  assign _03139_ = \bapg_rd.w_ptr_r [2] ? _03138_ : _03135_;
  assign _03140_ = \bapg_rd.w_ptr_r [3] ? _03139_ : _03132_;
  assign _03141_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [2] : \MSYNC_1r1w.synth.nz.mem[16] [2];
  assign _03142_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [2] : \MSYNC_1r1w.synth.nz.mem[18] [2];
  assign _03143_ = \bapg_rd.w_ptr_r [1] ? _03142_ : _03141_;
  assign _03144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [2] : \MSYNC_1r1w.synth.nz.mem[20] [2];
  assign _03145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [2] : \MSYNC_1r1w.synth.nz.mem[22] [2];
  assign _03146_ = \bapg_rd.w_ptr_r [1] ? _03145_ : _03144_;
  assign _03147_ = \bapg_rd.w_ptr_r [2] ? _03146_ : _03143_;
  assign _03148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [2] : \MSYNC_1r1w.synth.nz.mem[24] [2];
  assign _03149_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [2] : \MSYNC_1r1w.synth.nz.mem[26] [2];
  assign _03150_ = \bapg_rd.w_ptr_r [1] ? _03149_ : _03148_;
  assign _03151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [2] : \MSYNC_1r1w.synth.nz.mem[28] [2];
  assign _03152_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [2] : \MSYNC_1r1w.synth.nz.mem[30] [2];
  assign _03153_ = \bapg_rd.w_ptr_r [1] ? _03152_ : _03151_;
  assign _03154_ = \bapg_rd.w_ptr_r [2] ? _03153_ : _03150_;
  assign _03155_ = \bapg_rd.w_ptr_r [3] ? _03154_ : _03147_;
  assign _03156_ = \bapg_rd.w_ptr_r [4] ? _03155_ : _03140_;
  assign _03157_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [2] : \MSYNC_1r1w.synth.nz.mem[32] [2];
  assign _03158_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [2] : \MSYNC_1r1w.synth.nz.mem[34] [2];
  assign _03159_ = \bapg_rd.w_ptr_r [1] ? _03158_ : _03157_;
  assign _03160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [2] : \MSYNC_1r1w.synth.nz.mem[36] [2];
  assign _03161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [2] : \MSYNC_1r1w.synth.nz.mem[38] [2];
  assign _03162_ = \bapg_rd.w_ptr_r [1] ? _03161_ : _03160_;
  assign _03163_ = \bapg_rd.w_ptr_r [2] ? _03162_ : _03159_;
  assign _03164_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [2] : \MSYNC_1r1w.synth.nz.mem[40] [2];
  assign _03165_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [2] : \MSYNC_1r1w.synth.nz.mem[42] [2];
  assign _03166_ = \bapg_rd.w_ptr_r [1] ? _03165_ : _03164_;
  assign _03167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [2] : \MSYNC_1r1w.synth.nz.mem[44] [2];
  assign _03168_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [2] : \MSYNC_1r1w.synth.nz.mem[46] [2];
  assign _03169_ = \bapg_rd.w_ptr_r [1] ? _03168_ : _03167_;
  assign _03170_ = \bapg_rd.w_ptr_r [2] ? _03169_ : _03166_;
  assign _03171_ = \bapg_rd.w_ptr_r [3] ? _03170_ : _03163_;
  assign _03172_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [2] : \MSYNC_1r1w.synth.nz.mem[48] [2];
  assign _03173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [2] : \MSYNC_1r1w.synth.nz.mem[50] [2];
  assign _03174_ = \bapg_rd.w_ptr_r [1] ? _03173_ : _03172_;
  assign _03175_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [2] : \MSYNC_1r1w.synth.nz.mem[52] [2];
  assign _03176_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [2] : \MSYNC_1r1w.synth.nz.mem[54] [2];
  assign _03177_ = \bapg_rd.w_ptr_r [1] ? _03176_ : _03175_;
  assign _03178_ = \bapg_rd.w_ptr_r [2] ? _03177_ : _03174_;
  assign _03179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [2] : \MSYNC_1r1w.synth.nz.mem[56] [2];
  assign _03180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [2] : \MSYNC_1r1w.synth.nz.mem[58] [2];
  assign _03181_ = \bapg_rd.w_ptr_r [1] ? _03180_ : _03179_;
  assign _03182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [2] : \MSYNC_1r1w.synth.nz.mem[60] [2];
  assign _03183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [2] : \MSYNC_1r1w.synth.nz.mem[62] [2];
  assign _03184_ = \bapg_rd.w_ptr_r [1] ? _03183_ : _03182_;
  assign _03185_ = \bapg_rd.w_ptr_r [2] ? _03184_ : _03181_;
  assign _03186_ = \bapg_rd.w_ptr_r [3] ? _03185_ : _03178_;
  assign _03187_ = \bapg_rd.w_ptr_r [4] ? _03186_ : _03171_;
  assign _03188_ = \bapg_rd.w_ptr_r [5] ? _03187_ : _03156_;
  assign _03189_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [2] : \MSYNC_1r1w.synth.nz.mem[64] [2];
  assign _03190_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [2] : \MSYNC_1r1w.synth.nz.mem[66] [2];
  assign _03191_ = \bapg_rd.w_ptr_r [1] ? _03190_ : _03189_;
  assign _03192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [2] : \MSYNC_1r1w.synth.nz.mem[68] [2];
  assign _03193_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [2] : \MSYNC_1r1w.synth.nz.mem[70] [2];
  assign _03194_ = \bapg_rd.w_ptr_r [1] ? _03193_ : _03192_;
  assign _03195_ = \bapg_rd.w_ptr_r [2] ? _03194_ : _03191_;
  assign _03196_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [2] : \MSYNC_1r1w.synth.nz.mem[72] [2];
  assign _03197_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [2] : \MSYNC_1r1w.synth.nz.mem[74] [2];
  assign _03198_ = \bapg_rd.w_ptr_r [1] ? _03197_ : _03196_;
  assign _03199_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [2] : \MSYNC_1r1w.synth.nz.mem[76] [2];
  assign _03200_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [2] : \MSYNC_1r1w.synth.nz.mem[78] [2];
  assign _03201_ = \bapg_rd.w_ptr_r [1] ? _03200_ : _03199_;
  assign _03202_ = \bapg_rd.w_ptr_r [2] ? _03201_ : _03198_;
  assign _03203_ = \bapg_rd.w_ptr_r [3] ? _03202_ : _03195_;
  assign _03204_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [2] : \MSYNC_1r1w.synth.nz.mem[80] [2];
  assign _03205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [2] : \MSYNC_1r1w.synth.nz.mem[82] [2];
  assign _03206_ = \bapg_rd.w_ptr_r [1] ? _03205_ : _03204_;
  assign _03207_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [2] : \MSYNC_1r1w.synth.nz.mem[84] [2];
  assign _03208_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [2] : \MSYNC_1r1w.synth.nz.mem[86] [2];
  assign _03209_ = \bapg_rd.w_ptr_r [1] ? _03208_ : _03207_;
  assign _03210_ = \bapg_rd.w_ptr_r [2] ? _03209_ : _03206_;
  assign _03211_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [2] : \MSYNC_1r1w.synth.nz.mem[88] [2];
  assign _03212_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [2] : \MSYNC_1r1w.synth.nz.mem[90] [2];
  assign _03213_ = \bapg_rd.w_ptr_r [1] ? _03212_ : _03211_;
  assign _03214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [2] : \MSYNC_1r1w.synth.nz.mem[92] [2];
  assign _03215_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [2] : \MSYNC_1r1w.synth.nz.mem[94] [2];
  assign _03216_ = \bapg_rd.w_ptr_r [1] ? _03215_ : _03214_;
  assign _03217_ = \bapg_rd.w_ptr_r [2] ? _03216_ : _03213_;
  assign _03218_ = \bapg_rd.w_ptr_r [3] ? _03217_ : _03210_;
  assign _03219_ = \bapg_rd.w_ptr_r [4] ? _03218_ : _03203_;
  assign _03220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [2] : \MSYNC_1r1w.synth.nz.mem[96] [2];
  assign _03221_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [2] : \MSYNC_1r1w.synth.nz.mem[98] [2];
  assign _03222_ = \bapg_rd.w_ptr_r [1] ? _03221_ : _03220_;
  assign _03223_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [2] : \MSYNC_1r1w.synth.nz.mem[100] [2];
  assign _03224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [2] : \MSYNC_1r1w.synth.nz.mem[102] [2];
  assign _03225_ = \bapg_rd.w_ptr_r [1] ? _03224_ : _03223_;
  assign _03226_ = \bapg_rd.w_ptr_r [2] ? _03225_ : _03222_;
  assign _03227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [2] : \MSYNC_1r1w.synth.nz.mem[104] [2];
  assign _03228_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [2] : \MSYNC_1r1w.synth.nz.mem[106] [2];
  assign _03229_ = \bapg_rd.w_ptr_r [1] ? _03228_ : _03227_;
  assign _03230_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [2] : \MSYNC_1r1w.synth.nz.mem[108] [2];
  assign _03231_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [2] : \MSYNC_1r1w.synth.nz.mem[110] [2];
  assign _03232_ = \bapg_rd.w_ptr_r [1] ? _03231_ : _03230_;
  assign _03233_ = \bapg_rd.w_ptr_r [2] ? _03232_ : _03229_;
  assign _03234_ = \bapg_rd.w_ptr_r [3] ? _03233_ : _03226_;
  assign _03235_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [2] : \MSYNC_1r1w.synth.nz.mem[112] [2];
  assign _03236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [2] : \MSYNC_1r1w.synth.nz.mem[114] [2];
  assign _03237_ = \bapg_rd.w_ptr_r [1] ? _03236_ : _03235_;
  assign _03238_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [2] : \MSYNC_1r1w.synth.nz.mem[116] [2];
  assign _03239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [2] : \MSYNC_1r1w.synth.nz.mem[118] [2];
  assign _03240_ = \bapg_rd.w_ptr_r [1] ? _03239_ : _03238_;
  assign _03241_ = \bapg_rd.w_ptr_r [2] ? _03240_ : _03237_;
  assign _03242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [2] : \MSYNC_1r1w.synth.nz.mem[120] [2];
  assign _03243_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [2] : \MSYNC_1r1w.synth.nz.mem[122] [2];
  assign _03244_ = \bapg_rd.w_ptr_r [1] ? _03243_ : _03242_;
  assign _03245_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [2] : \MSYNC_1r1w.synth.nz.mem[124] [2];
  assign _03246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [2] : \MSYNC_1r1w.synth.nz.mem[126] [2];
  assign _03247_ = \bapg_rd.w_ptr_r [1] ? _03246_ : _03245_;
  assign _03248_ = \bapg_rd.w_ptr_r [2] ? _03247_ : _03244_;
  assign _03249_ = \bapg_rd.w_ptr_r [3] ? _03248_ : _03241_;
  assign _03250_ = \bapg_rd.w_ptr_r [4] ? _03249_ : _03234_;
  assign _03251_ = \bapg_rd.w_ptr_r [5] ? _03250_ : _03219_;
  assign _03252_ = \bapg_rd.w_ptr_r [6] ? _03251_ : _03188_;
  assign _03253_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [2] : \MSYNC_1r1w.synth.nz.mem[128] [2];
  assign _03254_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [2] : \MSYNC_1r1w.synth.nz.mem[130] [2];
  assign _03255_ = \bapg_rd.w_ptr_r [1] ? _03254_ : _03253_;
  assign _03256_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [2] : \MSYNC_1r1w.synth.nz.mem[132] [2];
  assign _03257_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [2] : \MSYNC_1r1w.synth.nz.mem[134] [2];
  assign _03258_ = \bapg_rd.w_ptr_r [1] ? _03257_ : _03256_;
  assign _03259_ = \bapg_rd.w_ptr_r [2] ? _03258_ : _03255_;
  assign _03260_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [2] : \MSYNC_1r1w.synth.nz.mem[136] [2];
  assign _03261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [2] : \MSYNC_1r1w.synth.nz.mem[138] [2];
  assign _03262_ = \bapg_rd.w_ptr_r [1] ? _03261_ : _03260_;
  assign _03263_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [2] : \MSYNC_1r1w.synth.nz.mem[140] [2];
  assign _03264_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [2] : \MSYNC_1r1w.synth.nz.mem[142] [2];
  assign _03265_ = \bapg_rd.w_ptr_r [1] ? _03264_ : _03263_;
  assign _03266_ = \bapg_rd.w_ptr_r [2] ? _03265_ : _03262_;
  assign _03267_ = \bapg_rd.w_ptr_r [3] ? _03266_ : _03259_;
  assign _03268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [2] : \MSYNC_1r1w.synth.nz.mem[144] [2];
  assign _03269_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [2] : \MSYNC_1r1w.synth.nz.mem[146] [2];
  assign _03270_ = \bapg_rd.w_ptr_r [1] ? _03269_ : _03268_;
  assign _03271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [2] : \MSYNC_1r1w.synth.nz.mem[148] [2];
  assign _03272_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [2] : \MSYNC_1r1w.synth.nz.mem[150] [2];
  assign _03273_ = \bapg_rd.w_ptr_r [1] ? _03272_ : _03271_;
  assign _03274_ = \bapg_rd.w_ptr_r [2] ? _03273_ : _03270_;
  assign _03275_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [2] : \MSYNC_1r1w.synth.nz.mem[152] [2];
  assign _03276_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [2] : \MSYNC_1r1w.synth.nz.mem[154] [2];
  assign _03277_ = \bapg_rd.w_ptr_r [1] ? _03276_ : _03275_;
  assign _03278_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [2] : \MSYNC_1r1w.synth.nz.mem[156] [2];
  assign _03279_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [2] : \MSYNC_1r1w.synth.nz.mem[158] [2];
  assign _03280_ = \bapg_rd.w_ptr_r [1] ? _03279_ : _03278_;
  assign _03281_ = \bapg_rd.w_ptr_r [2] ? _03280_ : _03277_;
  assign _03282_ = \bapg_rd.w_ptr_r [3] ? _03281_ : _03274_;
  assign _03283_ = \bapg_rd.w_ptr_r [4] ? _03282_ : _03267_;
  assign _03284_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [2] : \MSYNC_1r1w.synth.nz.mem[160] [2];
  assign _03285_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [2] : \MSYNC_1r1w.synth.nz.mem[162] [2];
  assign _03286_ = \bapg_rd.w_ptr_r [1] ? _03285_ : _03284_;
  assign _03287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [2] : \MSYNC_1r1w.synth.nz.mem[164] [2];
  assign _03288_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [2] : \MSYNC_1r1w.synth.nz.mem[166] [2];
  assign _03289_ = \bapg_rd.w_ptr_r [1] ? _03288_ : _03287_;
  assign _03290_ = \bapg_rd.w_ptr_r [2] ? _03289_ : _03286_;
  assign _03291_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [2] : \MSYNC_1r1w.synth.nz.mem[168] [2];
  assign _03292_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [2] : \MSYNC_1r1w.synth.nz.mem[170] [2];
  assign _03293_ = \bapg_rd.w_ptr_r [1] ? _03292_ : _03291_;
  assign _03294_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [2] : \MSYNC_1r1w.synth.nz.mem[172] [2];
  assign _03295_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [2] : \MSYNC_1r1w.synth.nz.mem[174] [2];
  assign _03296_ = \bapg_rd.w_ptr_r [1] ? _03295_ : _03294_;
  assign _03297_ = \bapg_rd.w_ptr_r [2] ? _03296_ : _03293_;
  assign _03298_ = \bapg_rd.w_ptr_r [3] ? _03297_ : _03290_;
  assign _03299_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [2] : \MSYNC_1r1w.synth.nz.mem[176] [2];
  assign _03300_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [2] : \MSYNC_1r1w.synth.nz.mem[178] [2];
  assign _03301_ = \bapg_rd.w_ptr_r [1] ? _03300_ : _03299_;
  assign _03302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [2] : \MSYNC_1r1w.synth.nz.mem[180] [2];
  assign _03303_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [2] : \MSYNC_1r1w.synth.nz.mem[182] [2];
  assign _03304_ = \bapg_rd.w_ptr_r [1] ? _03303_ : _03302_;
  assign _03305_ = \bapg_rd.w_ptr_r [2] ? _03304_ : _03301_;
  assign _03306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [2] : \MSYNC_1r1w.synth.nz.mem[184] [2];
  assign _03307_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [2] : \MSYNC_1r1w.synth.nz.mem[186] [2];
  assign _03308_ = \bapg_rd.w_ptr_r [1] ? _03307_ : _03306_;
  assign _03309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [2] : \MSYNC_1r1w.synth.nz.mem[188] [2];
  assign _03310_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [2] : \MSYNC_1r1w.synth.nz.mem[190] [2];
  assign _03311_ = \bapg_rd.w_ptr_r [1] ? _03310_ : _03309_;
  assign _03312_ = \bapg_rd.w_ptr_r [2] ? _03311_ : _03308_;
  assign _03313_ = \bapg_rd.w_ptr_r [3] ? _03312_ : _03305_;
  assign _03314_ = \bapg_rd.w_ptr_r [4] ? _03313_ : _03298_;
  assign _03315_ = \bapg_rd.w_ptr_r [5] ? _03314_ : _03283_;
  assign _03316_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [2] : \MSYNC_1r1w.synth.nz.mem[192] [2];
  assign _03317_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [2] : \MSYNC_1r1w.synth.nz.mem[194] [2];
  assign _03318_ = \bapg_rd.w_ptr_r [1] ? _03317_ : _03316_;
  assign _03319_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [2] : \MSYNC_1r1w.synth.nz.mem[196] [2];
  assign _03320_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [2] : \MSYNC_1r1w.synth.nz.mem[198] [2];
  assign _03321_ = \bapg_rd.w_ptr_r [1] ? _03320_ : _03319_;
  assign _03322_ = \bapg_rd.w_ptr_r [2] ? _03321_ : _03318_;
  assign _03323_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [2] : \MSYNC_1r1w.synth.nz.mem[200] [2];
  assign _03324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [2] : \MSYNC_1r1w.synth.nz.mem[202] [2];
  assign _03325_ = \bapg_rd.w_ptr_r [1] ? _03324_ : _03323_;
  assign _03326_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [2] : \MSYNC_1r1w.synth.nz.mem[204] [2];
  assign _03327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [2] : \MSYNC_1r1w.synth.nz.mem[206] [2];
  assign _03328_ = \bapg_rd.w_ptr_r [1] ? _03327_ : _03326_;
  assign _03329_ = \bapg_rd.w_ptr_r [2] ? _03328_ : _03325_;
  assign _03330_ = \bapg_rd.w_ptr_r [3] ? _03329_ : _03322_;
  assign _03331_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [2] : \MSYNC_1r1w.synth.nz.mem[208] [2];
  assign _03332_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [2] : \MSYNC_1r1w.synth.nz.mem[210] [2];
  assign _03333_ = \bapg_rd.w_ptr_r [1] ? _03332_ : _03331_;
  assign _03334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [2] : \MSYNC_1r1w.synth.nz.mem[212] [2];
  assign _03335_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [2] : \MSYNC_1r1w.synth.nz.mem[214] [2];
  assign _03336_ = \bapg_rd.w_ptr_r [1] ? _03335_ : _03334_;
  assign _03337_ = \bapg_rd.w_ptr_r [2] ? _03336_ : _03333_;
  assign _03338_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [2] : \MSYNC_1r1w.synth.nz.mem[216] [2];
  assign _03339_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [2] : \MSYNC_1r1w.synth.nz.mem[218] [2];
  assign _03340_ = \bapg_rd.w_ptr_r [1] ? _03339_ : _03338_;
  assign _03341_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [2] : \MSYNC_1r1w.synth.nz.mem[220] [2];
  assign _03342_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [2] : \MSYNC_1r1w.synth.nz.mem[222] [2];
  assign _03343_ = \bapg_rd.w_ptr_r [1] ? _03342_ : _03341_;
  assign _03344_ = \bapg_rd.w_ptr_r [2] ? _03343_ : _03340_;
  assign _03345_ = \bapg_rd.w_ptr_r [3] ? _03344_ : _03337_;
  assign _03346_ = \bapg_rd.w_ptr_r [4] ? _03345_ : _03330_;
  assign _03347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [2] : \MSYNC_1r1w.synth.nz.mem[224] [2];
  assign _03348_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [2] : \MSYNC_1r1w.synth.nz.mem[226] [2];
  assign _03349_ = \bapg_rd.w_ptr_r [1] ? _03348_ : _03347_;
  assign _03350_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [2] : \MSYNC_1r1w.synth.nz.mem[228] [2];
  assign _03351_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [2] : \MSYNC_1r1w.synth.nz.mem[230] [2];
  assign _03352_ = \bapg_rd.w_ptr_r [1] ? _03351_ : _03350_;
  assign _03353_ = \bapg_rd.w_ptr_r [2] ? _03352_ : _03349_;
  assign _03354_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [2] : \MSYNC_1r1w.synth.nz.mem[232] [2];
  assign _03355_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [2] : \MSYNC_1r1w.synth.nz.mem[234] [2];
  assign _03356_ = \bapg_rd.w_ptr_r [1] ? _03355_ : _03354_;
  assign _03357_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [2] : \MSYNC_1r1w.synth.nz.mem[236] [2];
  assign _03358_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [2] : \MSYNC_1r1w.synth.nz.mem[238] [2];
  assign _03359_ = \bapg_rd.w_ptr_r [1] ? _03358_ : _03357_;
  assign _03360_ = \bapg_rd.w_ptr_r [2] ? _03359_ : _03356_;
  assign _03361_ = \bapg_rd.w_ptr_r [3] ? _03360_ : _03353_;
  assign _03362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [2] : \MSYNC_1r1w.synth.nz.mem[240] [2];
  assign _03363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [2] : \MSYNC_1r1w.synth.nz.mem[242] [2];
  assign _03364_ = \bapg_rd.w_ptr_r [1] ? _03363_ : _03362_;
  assign _03365_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [2] : \MSYNC_1r1w.synth.nz.mem[244] [2];
  assign _03366_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [2] : \MSYNC_1r1w.synth.nz.mem[246] [2];
  assign _03367_ = \bapg_rd.w_ptr_r [1] ? _03366_ : _03365_;
  assign _03368_ = \bapg_rd.w_ptr_r [2] ? _03367_ : _03364_;
  assign _03369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [2] : \MSYNC_1r1w.synth.nz.mem[248] [2];
  assign _03370_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [2] : \MSYNC_1r1w.synth.nz.mem[250] [2];
  assign _03371_ = \bapg_rd.w_ptr_r [1] ? _03370_ : _03369_;
  assign _03372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [2] : \MSYNC_1r1w.synth.nz.mem[252] [2];
  assign _03373_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [2] : \MSYNC_1r1w.synth.nz.mem[254] [2];
  assign _03374_ = \bapg_rd.w_ptr_r [1] ? _03373_ : _03372_;
  assign _03375_ = \bapg_rd.w_ptr_r [2] ? _03374_ : _03371_;
  assign _03376_ = \bapg_rd.w_ptr_r [3] ? _03375_ : _03368_;
  assign _03377_ = \bapg_rd.w_ptr_r [4] ? _03376_ : _03361_;
  assign _03378_ = \bapg_rd.w_ptr_r [5] ? _03377_ : _03346_;
  assign _03379_ = \bapg_rd.w_ptr_r [6] ? _03378_ : _03315_;
  assign _03380_ = \bapg_rd.w_ptr_r [7] ? _03379_ : _03252_;
  assign _03381_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [2] : \MSYNC_1r1w.synth.nz.mem[256] [2];
  assign _03382_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [2] : \MSYNC_1r1w.synth.nz.mem[258] [2];
  assign _03383_ = \bapg_rd.w_ptr_r [1] ? _03382_ : _03381_;
  assign _03384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [2] : \MSYNC_1r1w.synth.nz.mem[260] [2];
  assign _03385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [2] : \MSYNC_1r1w.synth.nz.mem[262] [2];
  assign _03386_ = \bapg_rd.w_ptr_r [1] ? _03385_ : _03384_;
  assign _03387_ = \bapg_rd.w_ptr_r [2] ? _03386_ : _03383_;
  assign _03388_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [2] : \MSYNC_1r1w.synth.nz.mem[264] [2];
  assign _03389_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [2] : \MSYNC_1r1w.synth.nz.mem[266] [2];
  assign _03390_ = \bapg_rd.w_ptr_r [1] ? _03389_ : _03388_;
  assign _03391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [2] : \MSYNC_1r1w.synth.nz.mem[268] [2];
  assign _03392_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [2] : \MSYNC_1r1w.synth.nz.mem[270] [2];
  assign _03393_ = \bapg_rd.w_ptr_r [1] ? _03392_ : _03391_;
  assign _03394_ = \bapg_rd.w_ptr_r [2] ? _03393_ : _03390_;
  assign _03395_ = \bapg_rd.w_ptr_r [3] ? _03394_ : _03387_;
  assign _03396_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [2] : \MSYNC_1r1w.synth.nz.mem[272] [2];
  assign _03397_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [2] : \MSYNC_1r1w.synth.nz.mem[274] [2];
  assign _03398_ = \bapg_rd.w_ptr_r [1] ? _03397_ : _03396_;
  assign _03399_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [2] : \MSYNC_1r1w.synth.nz.mem[276] [2];
  assign _03400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [2] : \MSYNC_1r1w.synth.nz.mem[278] [2];
  assign _03401_ = \bapg_rd.w_ptr_r [1] ? _03400_ : _03399_;
  assign _03402_ = \bapg_rd.w_ptr_r [2] ? _03401_ : _03398_;
  assign _03403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [2] : \MSYNC_1r1w.synth.nz.mem[280] [2];
  assign _03404_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [2] : \MSYNC_1r1w.synth.nz.mem[282] [2];
  assign _03405_ = \bapg_rd.w_ptr_r [1] ? _03404_ : _03403_;
  assign _03406_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [2] : \MSYNC_1r1w.synth.nz.mem[284] [2];
  assign _03407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [2] : \MSYNC_1r1w.synth.nz.mem[286] [2];
  assign _03408_ = \bapg_rd.w_ptr_r [1] ? _03407_ : _03406_;
  assign _03409_ = \bapg_rd.w_ptr_r [2] ? _03408_ : _03405_;
  assign _03410_ = \bapg_rd.w_ptr_r [3] ? _03409_ : _03402_;
  assign _03411_ = \bapg_rd.w_ptr_r [4] ? _03410_ : _03395_;
  assign _03412_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [2] : \MSYNC_1r1w.synth.nz.mem[288] [2];
  assign _03413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [2] : \MSYNC_1r1w.synth.nz.mem[290] [2];
  assign _03414_ = \bapg_rd.w_ptr_r [1] ? _03413_ : _03412_;
  assign _03415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [2] : \MSYNC_1r1w.synth.nz.mem[292] [2];
  assign _03416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [2] : \MSYNC_1r1w.synth.nz.mem[294] [2];
  assign _03417_ = \bapg_rd.w_ptr_r [1] ? _03416_ : _03415_;
  assign _03418_ = \bapg_rd.w_ptr_r [2] ? _03417_ : _03414_;
  assign _03419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [2] : \MSYNC_1r1w.synth.nz.mem[296] [2];
  assign _03420_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [2] : \MSYNC_1r1w.synth.nz.mem[298] [2];
  assign _03421_ = \bapg_rd.w_ptr_r [1] ? _03420_ : _03419_;
  assign _03422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [2] : \MSYNC_1r1w.synth.nz.mem[300] [2];
  assign _03423_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [2] : \MSYNC_1r1w.synth.nz.mem[302] [2];
  assign _03424_ = \bapg_rd.w_ptr_r [1] ? _03423_ : _03422_;
  assign _03425_ = \bapg_rd.w_ptr_r [2] ? _03424_ : _03421_;
  assign _03426_ = \bapg_rd.w_ptr_r [3] ? _03425_ : _03418_;
  assign _03427_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [2] : \MSYNC_1r1w.synth.nz.mem[304] [2];
  assign _03428_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [2] : \MSYNC_1r1w.synth.nz.mem[306] [2];
  assign _03429_ = \bapg_rd.w_ptr_r [1] ? _03428_ : _03427_;
  assign _03430_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [2] : \MSYNC_1r1w.synth.nz.mem[308] [2];
  assign _03431_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [2] : \MSYNC_1r1w.synth.nz.mem[310] [2];
  assign _03432_ = \bapg_rd.w_ptr_r [1] ? _03431_ : _03430_;
  assign _03433_ = \bapg_rd.w_ptr_r [2] ? _03432_ : _03429_;
  assign _03434_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [2] : \MSYNC_1r1w.synth.nz.mem[312] [2];
  assign _03435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [2] : \MSYNC_1r1w.synth.nz.mem[314] [2];
  assign _03436_ = \bapg_rd.w_ptr_r [1] ? _03435_ : _03434_;
  assign _03437_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [2] : \MSYNC_1r1w.synth.nz.mem[316] [2];
  assign _03438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [2] : \MSYNC_1r1w.synth.nz.mem[318] [2];
  assign _03439_ = \bapg_rd.w_ptr_r [1] ? _03438_ : _03437_;
  assign _03440_ = \bapg_rd.w_ptr_r [2] ? _03439_ : _03436_;
  assign _03441_ = \bapg_rd.w_ptr_r [3] ? _03440_ : _03433_;
  assign _03442_ = \bapg_rd.w_ptr_r [4] ? _03441_ : _03426_;
  assign _03443_ = \bapg_rd.w_ptr_r [5] ? _03442_ : _03411_;
  assign _03444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [2] : \MSYNC_1r1w.synth.nz.mem[320] [2];
  assign _03445_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [2] : \MSYNC_1r1w.synth.nz.mem[322] [2];
  assign _03446_ = \bapg_rd.w_ptr_r [1] ? _03445_ : _03444_;
  assign _03447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [2] : \MSYNC_1r1w.synth.nz.mem[324] [2];
  assign _03448_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [2] : \MSYNC_1r1w.synth.nz.mem[326] [2];
  assign _03449_ = \bapg_rd.w_ptr_r [1] ? _03448_ : _03447_;
  assign _03450_ = \bapg_rd.w_ptr_r [2] ? _03449_ : _03446_;
  assign _03451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [2] : \MSYNC_1r1w.synth.nz.mem[328] [2];
  assign _03452_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [2] : \MSYNC_1r1w.synth.nz.mem[330] [2];
  assign _03453_ = \bapg_rd.w_ptr_r [1] ? _03452_ : _03451_;
  assign _03454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [2] : \MSYNC_1r1w.synth.nz.mem[332] [2];
  assign _03455_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [2] : \MSYNC_1r1w.synth.nz.mem[334] [2];
  assign _03456_ = \bapg_rd.w_ptr_r [1] ? _03455_ : _03454_;
  assign _03457_ = \bapg_rd.w_ptr_r [2] ? _03456_ : _03453_;
  assign _03458_ = \bapg_rd.w_ptr_r [3] ? _03457_ : _03450_;
  assign _03459_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [2] : \MSYNC_1r1w.synth.nz.mem[336] [2];
  assign _03460_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [2] : \MSYNC_1r1w.synth.nz.mem[338] [2];
  assign _03461_ = \bapg_rd.w_ptr_r [1] ? _03460_ : _03459_;
  assign _03462_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [2] : \MSYNC_1r1w.synth.nz.mem[340] [2];
  assign _03463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [2] : \MSYNC_1r1w.synth.nz.mem[342] [2];
  assign _03464_ = \bapg_rd.w_ptr_r [1] ? _03463_ : _03462_;
  assign _03465_ = \bapg_rd.w_ptr_r [2] ? _03464_ : _03461_;
  assign _03466_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [2] : \MSYNC_1r1w.synth.nz.mem[344] [2];
  assign _03467_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [2] : \MSYNC_1r1w.synth.nz.mem[346] [2];
  assign _03468_ = \bapg_rd.w_ptr_r [1] ? _03467_ : _03466_;
  assign _03469_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [2] : \MSYNC_1r1w.synth.nz.mem[348] [2];
  assign _03470_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [2] : \MSYNC_1r1w.synth.nz.mem[350] [2];
  assign _03471_ = \bapg_rd.w_ptr_r [1] ? _03470_ : _03469_;
  assign _03472_ = \bapg_rd.w_ptr_r [2] ? _03471_ : _03468_;
  assign _03473_ = \bapg_rd.w_ptr_r [3] ? _03472_ : _03465_;
  assign _03474_ = \bapg_rd.w_ptr_r [4] ? _03473_ : _03458_;
  assign _03475_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [2] : \MSYNC_1r1w.synth.nz.mem[352] [2];
  assign _03476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [2] : \MSYNC_1r1w.synth.nz.mem[354] [2];
  assign _03477_ = \bapg_rd.w_ptr_r [1] ? _03476_ : _03475_;
  assign _03478_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [2] : \MSYNC_1r1w.synth.nz.mem[356] [2];
  assign _03479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [2] : \MSYNC_1r1w.synth.nz.mem[358] [2];
  assign _03480_ = \bapg_rd.w_ptr_r [1] ? _03479_ : _03478_;
  assign _03481_ = \bapg_rd.w_ptr_r [2] ? _03480_ : _03477_;
  assign _03482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [2] : \MSYNC_1r1w.synth.nz.mem[360] [2];
  assign _03483_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [2] : \MSYNC_1r1w.synth.nz.mem[362] [2];
  assign _03484_ = \bapg_rd.w_ptr_r [1] ? _03483_ : _03482_;
  assign _03485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [2] : \MSYNC_1r1w.synth.nz.mem[364] [2];
  assign _03486_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [2] : \MSYNC_1r1w.synth.nz.mem[366] [2];
  assign _03487_ = \bapg_rd.w_ptr_r [1] ? _03486_ : _03485_;
  assign _03488_ = \bapg_rd.w_ptr_r [2] ? _03487_ : _03484_;
  assign _03489_ = \bapg_rd.w_ptr_r [3] ? _03488_ : _03481_;
  assign _03490_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [2] : \MSYNC_1r1w.synth.nz.mem[368] [2];
  assign _03491_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [2] : \MSYNC_1r1w.synth.nz.mem[370] [2];
  assign _03492_ = \bapg_rd.w_ptr_r [1] ? _03491_ : _03490_;
  assign _03493_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [2] : \MSYNC_1r1w.synth.nz.mem[372] [2];
  assign _03494_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [2] : \MSYNC_1r1w.synth.nz.mem[374] [2];
  assign _03495_ = \bapg_rd.w_ptr_r [1] ? _03494_ : _03493_;
  assign _03496_ = \bapg_rd.w_ptr_r [2] ? _03495_ : _03492_;
  assign _03497_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [2] : \MSYNC_1r1w.synth.nz.mem[376] [2];
  assign _03498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [2] : \MSYNC_1r1w.synth.nz.mem[378] [2];
  assign _03499_ = \bapg_rd.w_ptr_r [1] ? _03498_ : _03497_;
  assign _03500_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [2] : \MSYNC_1r1w.synth.nz.mem[380] [2];
  assign _03501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [2] : \MSYNC_1r1w.synth.nz.mem[382] [2];
  assign _03502_ = \bapg_rd.w_ptr_r [1] ? _03501_ : _03500_;
  assign _03503_ = \bapg_rd.w_ptr_r [2] ? _03502_ : _03499_;
  assign _03504_ = \bapg_rd.w_ptr_r [3] ? _03503_ : _03496_;
  assign _03505_ = \bapg_rd.w_ptr_r [4] ? _03504_ : _03489_;
  assign _03506_ = \bapg_rd.w_ptr_r [5] ? _03505_ : _03474_;
  assign _03507_ = \bapg_rd.w_ptr_r [6] ? _03506_ : _03443_;
  assign _03508_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [2] : \MSYNC_1r1w.synth.nz.mem[384] [2];
  assign _03509_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [2] : \MSYNC_1r1w.synth.nz.mem[386] [2];
  assign _03510_ = \bapg_rd.w_ptr_r [1] ? _03509_ : _03508_;
  assign _03511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [2] : \MSYNC_1r1w.synth.nz.mem[388] [2];
  assign _03512_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [2] : \MSYNC_1r1w.synth.nz.mem[390] [2];
  assign _03513_ = \bapg_rd.w_ptr_r [1] ? _03512_ : _03511_;
  assign _03514_ = \bapg_rd.w_ptr_r [2] ? _03513_ : _03510_;
  assign _03515_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [2] : \MSYNC_1r1w.synth.nz.mem[392] [2];
  assign _03516_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [2] : \MSYNC_1r1w.synth.nz.mem[394] [2];
  assign _03517_ = \bapg_rd.w_ptr_r [1] ? _03516_ : _03515_;
  assign _03518_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [2] : \MSYNC_1r1w.synth.nz.mem[396] [2];
  assign _03519_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [2] : \MSYNC_1r1w.synth.nz.mem[398] [2];
  assign _03520_ = \bapg_rd.w_ptr_r [1] ? _03519_ : _03518_;
  assign _03521_ = \bapg_rd.w_ptr_r [2] ? _03520_ : _03517_;
  assign _03522_ = \bapg_rd.w_ptr_r [3] ? _03521_ : _03514_;
  assign _03523_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [2] : \MSYNC_1r1w.synth.nz.mem[400] [2];
  assign _03524_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [2] : \MSYNC_1r1w.synth.nz.mem[402] [2];
  assign _03525_ = \bapg_rd.w_ptr_r [1] ? _03524_ : _03523_;
  assign _03526_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [2] : \MSYNC_1r1w.synth.nz.mem[404] [2];
  assign _03527_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [2] : \MSYNC_1r1w.synth.nz.mem[406] [2];
  assign _03528_ = \bapg_rd.w_ptr_r [1] ? _03527_ : _03526_;
  assign _03529_ = \bapg_rd.w_ptr_r [2] ? _03528_ : _03525_;
  assign _03530_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [2] : \MSYNC_1r1w.synth.nz.mem[408] [2];
  assign _03531_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [2] : \MSYNC_1r1w.synth.nz.mem[410] [2];
  assign _03532_ = \bapg_rd.w_ptr_r [1] ? _03531_ : _03530_;
  assign _03533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [2] : \MSYNC_1r1w.synth.nz.mem[412] [2];
  assign _03534_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [2] : \MSYNC_1r1w.synth.nz.mem[414] [2];
  assign _03535_ = \bapg_rd.w_ptr_r [1] ? _03534_ : _03533_;
  assign _03536_ = \bapg_rd.w_ptr_r [2] ? _03535_ : _03532_;
  assign _03537_ = \bapg_rd.w_ptr_r [3] ? _03536_ : _03529_;
  assign _03538_ = \bapg_rd.w_ptr_r [4] ? _03537_ : _03522_;
  assign _03539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [2] : \MSYNC_1r1w.synth.nz.mem[416] [2];
  assign _03540_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [2] : \MSYNC_1r1w.synth.nz.mem[418] [2];
  assign _03541_ = \bapg_rd.w_ptr_r [1] ? _03540_ : _03539_;
  assign _03542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [2] : \MSYNC_1r1w.synth.nz.mem[420] [2];
  assign _03543_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [2] : \MSYNC_1r1w.synth.nz.mem[422] [2];
  assign _03544_ = \bapg_rd.w_ptr_r [1] ? _03543_ : _03542_;
  assign _03545_ = \bapg_rd.w_ptr_r [2] ? _03544_ : _03541_;
  assign _03546_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [2] : \MSYNC_1r1w.synth.nz.mem[424] [2];
  assign _03547_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [2] : \MSYNC_1r1w.synth.nz.mem[426] [2];
  assign _03548_ = \bapg_rd.w_ptr_r [1] ? _03547_ : _03546_;
  assign _03549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [2] : \MSYNC_1r1w.synth.nz.mem[428] [2];
  assign _03550_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [2] : \MSYNC_1r1w.synth.nz.mem[430] [2];
  assign _03551_ = \bapg_rd.w_ptr_r [1] ? _03550_ : _03549_;
  assign _03552_ = \bapg_rd.w_ptr_r [2] ? _03551_ : _03548_;
  assign _03553_ = \bapg_rd.w_ptr_r [3] ? _03552_ : _03545_;
  assign _03554_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [2] : \MSYNC_1r1w.synth.nz.mem[432] [2];
  assign _03555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [2] : \MSYNC_1r1w.synth.nz.mem[434] [2];
  assign _03556_ = \bapg_rd.w_ptr_r [1] ? _03555_ : _03554_;
  assign _03557_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [2] : \MSYNC_1r1w.synth.nz.mem[436] [2];
  assign _03558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [2] : \MSYNC_1r1w.synth.nz.mem[438] [2];
  assign _03559_ = \bapg_rd.w_ptr_r [1] ? _03558_ : _03557_;
  assign _03560_ = \bapg_rd.w_ptr_r [2] ? _03559_ : _03556_;
  assign _03561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [2] : \MSYNC_1r1w.synth.nz.mem[440] [2];
  assign _03562_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [2] : \MSYNC_1r1w.synth.nz.mem[442] [2];
  assign _03563_ = \bapg_rd.w_ptr_r [1] ? _03562_ : _03561_;
  assign _03564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [2] : \MSYNC_1r1w.synth.nz.mem[444] [2];
  assign _03565_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [2] : \MSYNC_1r1w.synth.nz.mem[446] [2];
  assign _03566_ = \bapg_rd.w_ptr_r [1] ? _03565_ : _03564_;
  assign _03567_ = \bapg_rd.w_ptr_r [2] ? _03566_ : _03563_;
  assign _03568_ = \bapg_rd.w_ptr_r [3] ? _03567_ : _03560_;
  assign _03569_ = \bapg_rd.w_ptr_r [4] ? _03568_ : _03553_;
  assign _03570_ = \bapg_rd.w_ptr_r [5] ? _03569_ : _03538_;
  assign _03571_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [2] : \MSYNC_1r1w.synth.nz.mem[448] [2];
  assign _03572_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [2] : \MSYNC_1r1w.synth.nz.mem[450] [2];
  assign _03573_ = \bapg_rd.w_ptr_r [1] ? _03572_ : _03571_;
  assign _03574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [2] : \MSYNC_1r1w.synth.nz.mem[452] [2];
  assign _03575_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [2] : \MSYNC_1r1w.synth.nz.mem[454] [2];
  assign _03576_ = \bapg_rd.w_ptr_r [1] ? _03575_ : _03574_;
  assign _03577_ = \bapg_rd.w_ptr_r [2] ? _03576_ : _03573_;
  assign _03578_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [2] : \MSYNC_1r1w.synth.nz.mem[456] [2];
  assign _03579_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [2] : \MSYNC_1r1w.synth.nz.mem[458] [2];
  assign _03580_ = \bapg_rd.w_ptr_r [1] ? _03579_ : _03578_;
  assign _03581_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [2] : \MSYNC_1r1w.synth.nz.mem[460] [2];
  assign _03582_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [2] : \MSYNC_1r1w.synth.nz.mem[462] [2];
  assign _03583_ = \bapg_rd.w_ptr_r [1] ? _03582_ : _03581_;
  assign _03584_ = \bapg_rd.w_ptr_r [2] ? _03583_ : _03580_;
  assign _03585_ = \bapg_rd.w_ptr_r [3] ? _03584_ : _03577_;
  assign _03586_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [2] : \MSYNC_1r1w.synth.nz.mem[464] [2];
  assign _03587_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [2] : \MSYNC_1r1w.synth.nz.mem[466] [2];
  assign _03588_ = \bapg_rd.w_ptr_r [1] ? _03587_ : _03586_;
  assign _03589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [2] : \MSYNC_1r1w.synth.nz.mem[468] [2];
  assign _03590_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [2] : \MSYNC_1r1w.synth.nz.mem[470] [2];
  assign _03591_ = \bapg_rd.w_ptr_r [1] ? _03590_ : _03589_;
  assign _03592_ = \bapg_rd.w_ptr_r [2] ? _03591_ : _03588_;
  assign _03593_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [2] : \MSYNC_1r1w.synth.nz.mem[472] [2];
  assign _03594_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [2] : \MSYNC_1r1w.synth.nz.mem[474] [2];
  assign _03595_ = \bapg_rd.w_ptr_r [1] ? _03594_ : _03593_;
  assign _03596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [2] : \MSYNC_1r1w.synth.nz.mem[476] [2];
  assign _03597_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [2] : \MSYNC_1r1w.synth.nz.mem[478] [2];
  assign _03598_ = \bapg_rd.w_ptr_r [1] ? _03597_ : _03596_;
  assign _03599_ = \bapg_rd.w_ptr_r [2] ? _03598_ : _03595_;
  assign _03600_ = \bapg_rd.w_ptr_r [3] ? _03599_ : _03592_;
  assign _03601_ = \bapg_rd.w_ptr_r [4] ? _03600_ : _03585_;
  assign _03602_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [2] : \MSYNC_1r1w.synth.nz.mem[480] [2];
  assign _03603_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [2] : \MSYNC_1r1w.synth.nz.mem[482] [2];
  assign _03604_ = \bapg_rd.w_ptr_r [1] ? _03603_ : _03602_;
  assign _03605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [2] : \MSYNC_1r1w.synth.nz.mem[484] [2];
  assign _03606_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [2] : \MSYNC_1r1w.synth.nz.mem[486] [2];
  assign _03607_ = \bapg_rd.w_ptr_r [1] ? _03606_ : _03605_;
  assign _03608_ = \bapg_rd.w_ptr_r [2] ? _03607_ : _03604_;
  assign _03609_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [2] : \MSYNC_1r1w.synth.nz.mem[488] [2];
  assign _03610_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [2] : \MSYNC_1r1w.synth.nz.mem[490] [2];
  assign _03611_ = \bapg_rd.w_ptr_r [1] ? _03610_ : _03609_;
  assign _03612_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [2] : \MSYNC_1r1w.synth.nz.mem[492] [2];
  assign _03613_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [2] : \MSYNC_1r1w.synth.nz.mem[494] [2];
  assign _03614_ = \bapg_rd.w_ptr_r [1] ? _03613_ : _03612_;
  assign _03615_ = \bapg_rd.w_ptr_r [2] ? _03614_ : _03611_;
  assign _03616_ = \bapg_rd.w_ptr_r [3] ? _03615_ : _03608_;
  assign _03617_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [2] : \MSYNC_1r1w.synth.nz.mem[496] [2];
  assign _03618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [2] : \MSYNC_1r1w.synth.nz.mem[498] [2];
  assign _03619_ = \bapg_rd.w_ptr_r [1] ? _03618_ : _03617_;
  assign _03620_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [2] : \MSYNC_1r1w.synth.nz.mem[500] [2];
  assign _03621_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [2] : \MSYNC_1r1w.synth.nz.mem[502] [2];
  assign _03622_ = \bapg_rd.w_ptr_r [1] ? _03621_ : _03620_;
  assign _03623_ = \bapg_rd.w_ptr_r [2] ? _03622_ : _03619_;
  assign _03624_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [2] : \MSYNC_1r1w.synth.nz.mem[504] [2];
  assign _03625_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [2] : \MSYNC_1r1w.synth.nz.mem[506] [2];
  assign _03626_ = \bapg_rd.w_ptr_r [1] ? _03625_ : _03624_;
  assign _03627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [2] : \MSYNC_1r1w.synth.nz.mem[508] [2];
  assign _03628_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [2] : \MSYNC_1r1w.synth.nz.mem[510] [2];
  assign _03629_ = \bapg_rd.w_ptr_r [1] ? _03628_ : _03627_;
  assign _03630_ = \bapg_rd.w_ptr_r [2] ? _03629_ : _03626_;
  assign _03631_ = \bapg_rd.w_ptr_r [3] ? _03630_ : _03623_;
  assign _03632_ = \bapg_rd.w_ptr_r [4] ? _03631_ : _03616_;
  assign _03633_ = \bapg_rd.w_ptr_r [5] ? _03632_ : _03601_;
  assign _03634_ = \bapg_rd.w_ptr_r [6] ? _03633_ : _03570_;
  assign _03635_ = \bapg_rd.w_ptr_r [7] ? _03634_ : _03507_;
  assign _03636_ = \bapg_rd.w_ptr_r [8] ? _03635_ : _03380_;
  assign _03637_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [2] : \MSYNC_1r1w.synth.nz.mem[512] [2];
  assign _03638_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [2] : \MSYNC_1r1w.synth.nz.mem[514] [2];
  assign _03639_ = \bapg_rd.w_ptr_r [1] ? _03638_ : _03637_;
  assign _03640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [2] : \MSYNC_1r1w.synth.nz.mem[516] [2];
  assign _03641_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [2] : \MSYNC_1r1w.synth.nz.mem[518] [2];
  assign _03642_ = \bapg_rd.w_ptr_r [1] ? _03641_ : _03640_;
  assign _03643_ = \bapg_rd.w_ptr_r [2] ? _03642_ : _03639_;
  assign _03644_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [2] : \MSYNC_1r1w.synth.nz.mem[520] [2];
  assign _03645_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [2] : \MSYNC_1r1w.synth.nz.mem[522] [2];
  assign _03646_ = \bapg_rd.w_ptr_r [1] ? _03645_ : _03644_;
  assign _03647_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [2] : \MSYNC_1r1w.synth.nz.mem[524] [2];
  assign _03648_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [2] : \MSYNC_1r1w.synth.nz.mem[526] [2];
  assign _03649_ = \bapg_rd.w_ptr_r [1] ? _03648_ : _03647_;
  assign _03650_ = \bapg_rd.w_ptr_r [2] ? _03649_ : _03646_;
  assign _03651_ = \bapg_rd.w_ptr_r [3] ? _03650_ : _03643_;
  assign _03652_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [2] : \MSYNC_1r1w.synth.nz.mem[528] [2];
  assign _03653_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [2] : \MSYNC_1r1w.synth.nz.mem[530] [2];
  assign _03654_ = \bapg_rd.w_ptr_r [1] ? _03653_ : _03652_;
  assign _03655_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [2] : \MSYNC_1r1w.synth.nz.mem[532] [2];
  assign _03656_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [2] : \MSYNC_1r1w.synth.nz.mem[534] [2];
  assign _03657_ = \bapg_rd.w_ptr_r [1] ? _03656_ : _03655_;
  assign _03658_ = \bapg_rd.w_ptr_r [2] ? _03657_ : _03654_;
  assign _03659_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [2] : \MSYNC_1r1w.synth.nz.mem[536] [2];
  assign _03660_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [2] : \MSYNC_1r1w.synth.nz.mem[538] [2];
  assign _03661_ = \bapg_rd.w_ptr_r [1] ? _03660_ : _03659_;
  assign _03662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [2] : \MSYNC_1r1w.synth.nz.mem[540] [2];
  assign _03663_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [2] : \MSYNC_1r1w.synth.nz.mem[542] [2];
  assign _03664_ = \bapg_rd.w_ptr_r [1] ? _03663_ : _03662_;
  assign _03665_ = \bapg_rd.w_ptr_r [2] ? _03664_ : _03661_;
  assign _03666_ = \bapg_rd.w_ptr_r [3] ? _03665_ : _03658_;
  assign _03667_ = \bapg_rd.w_ptr_r [4] ? _03666_ : _03651_;
  assign _03668_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [2] : \MSYNC_1r1w.synth.nz.mem[544] [2];
  assign _03669_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [2] : \MSYNC_1r1w.synth.nz.mem[546] [2];
  assign _03670_ = \bapg_rd.w_ptr_r [1] ? _03669_ : _03668_;
  assign _03671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [2] : \MSYNC_1r1w.synth.nz.mem[548] [2];
  assign _03672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [2] : \MSYNC_1r1w.synth.nz.mem[550] [2];
  assign _03673_ = \bapg_rd.w_ptr_r [1] ? _03672_ : _03671_;
  assign _03674_ = \bapg_rd.w_ptr_r [2] ? _03673_ : _03670_;
  assign _03675_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [2] : \MSYNC_1r1w.synth.nz.mem[552] [2];
  assign _03676_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [2] : \MSYNC_1r1w.synth.nz.mem[554] [2];
  assign _03677_ = \bapg_rd.w_ptr_r [1] ? _03676_ : _03675_;
  assign _03678_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [2] : \MSYNC_1r1w.synth.nz.mem[556] [2];
  assign _03679_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [2] : \MSYNC_1r1w.synth.nz.mem[558] [2];
  assign _03680_ = \bapg_rd.w_ptr_r [1] ? _03679_ : _03678_;
  assign _03681_ = \bapg_rd.w_ptr_r [2] ? _03680_ : _03677_;
  assign _03682_ = \bapg_rd.w_ptr_r [3] ? _03681_ : _03674_;
  assign _03683_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [2] : \MSYNC_1r1w.synth.nz.mem[560] [2];
  assign _03684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [2] : \MSYNC_1r1w.synth.nz.mem[562] [2];
  assign _03685_ = \bapg_rd.w_ptr_r [1] ? _03684_ : _03683_;
  assign _03686_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [2] : \MSYNC_1r1w.synth.nz.mem[564] [2];
  assign _03687_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [2] : \MSYNC_1r1w.synth.nz.mem[566] [2];
  assign _03688_ = \bapg_rd.w_ptr_r [1] ? _03687_ : _03686_;
  assign _03689_ = \bapg_rd.w_ptr_r [2] ? _03688_ : _03685_;
  assign _03690_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [2] : \MSYNC_1r1w.synth.nz.mem[568] [2];
  assign _03691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [2] : \MSYNC_1r1w.synth.nz.mem[570] [2];
  assign _03692_ = \bapg_rd.w_ptr_r [1] ? _03691_ : _03690_;
  assign _03693_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [2] : \MSYNC_1r1w.synth.nz.mem[572] [2];
  assign _03694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [2] : \MSYNC_1r1w.synth.nz.mem[574] [2];
  assign _03695_ = \bapg_rd.w_ptr_r [1] ? _03694_ : _03693_;
  assign _03696_ = \bapg_rd.w_ptr_r [2] ? _03695_ : _03692_;
  assign _03697_ = \bapg_rd.w_ptr_r [3] ? _03696_ : _03689_;
  assign _03698_ = \bapg_rd.w_ptr_r [4] ? _03697_ : _03682_;
  assign _03699_ = \bapg_rd.w_ptr_r [5] ? _03698_ : _03667_;
  assign _03700_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [2] : \MSYNC_1r1w.synth.nz.mem[576] [2];
  assign _03701_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [2] : \MSYNC_1r1w.synth.nz.mem[578] [2];
  assign _03702_ = \bapg_rd.w_ptr_r [1] ? _03701_ : _03700_;
  assign _03703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [2] : \MSYNC_1r1w.synth.nz.mem[580] [2];
  assign _03704_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [2] : \MSYNC_1r1w.synth.nz.mem[582] [2];
  assign _03705_ = \bapg_rd.w_ptr_r [1] ? _03704_ : _03703_;
  assign _03706_ = \bapg_rd.w_ptr_r [2] ? _03705_ : _03702_;
  assign _03707_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [2] : \MSYNC_1r1w.synth.nz.mem[584] [2];
  assign _03708_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [2] : \MSYNC_1r1w.synth.nz.mem[586] [2];
  assign _03709_ = \bapg_rd.w_ptr_r [1] ? _03708_ : _03707_;
  assign _03710_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [2] : \MSYNC_1r1w.synth.nz.mem[588] [2];
  assign _03711_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [2] : \MSYNC_1r1w.synth.nz.mem[590] [2];
  assign _03712_ = \bapg_rd.w_ptr_r [1] ? _03711_ : _03710_;
  assign _03713_ = \bapg_rd.w_ptr_r [2] ? _03712_ : _03709_;
  assign _03714_ = \bapg_rd.w_ptr_r [3] ? _03713_ : _03706_;
  assign _03715_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [2] : \MSYNC_1r1w.synth.nz.mem[592] [2];
  assign _03716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [2] : \MSYNC_1r1w.synth.nz.mem[594] [2];
  assign _03717_ = \bapg_rd.w_ptr_r [1] ? _03716_ : _03715_;
  assign _03718_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [2] : \MSYNC_1r1w.synth.nz.mem[596] [2];
  assign _03719_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [2] : \MSYNC_1r1w.synth.nz.mem[598] [2];
  assign _03720_ = \bapg_rd.w_ptr_r [1] ? _03719_ : _03718_;
  assign _03721_ = \bapg_rd.w_ptr_r [2] ? _03720_ : _03717_;
  assign _03722_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [2] : \MSYNC_1r1w.synth.nz.mem[600] [2];
  assign _03723_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [2] : \MSYNC_1r1w.synth.nz.mem[602] [2];
  assign _03724_ = \bapg_rd.w_ptr_r [1] ? _03723_ : _03722_;
  assign _03725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [2] : \MSYNC_1r1w.synth.nz.mem[604] [2];
  assign _03726_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [2] : \MSYNC_1r1w.synth.nz.mem[606] [2];
  assign _03727_ = \bapg_rd.w_ptr_r [1] ? _03726_ : _03725_;
  assign _03728_ = \bapg_rd.w_ptr_r [2] ? _03727_ : _03724_;
  assign _03729_ = \bapg_rd.w_ptr_r [3] ? _03728_ : _03721_;
  assign _03730_ = \bapg_rd.w_ptr_r [4] ? _03729_ : _03714_;
  assign _03731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [2] : \MSYNC_1r1w.synth.nz.mem[608] [2];
  assign _03732_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [2] : \MSYNC_1r1w.synth.nz.mem[610] [2];
  assign _03733_ = \bapg_rd.w_ptr_r [1] ? _03732_ : _03731_;
  assign _03734_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [2] : \MSYNC_1r1w.synth.nz.mem[612] [2];
  assign _03735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [2] : \MSYNC_1r1w.synth.nz.mem[614] [2];
  assign _03736_ = \bapg_rd.w_ptr_r [1] ? _03735_ : _03734_;
  assign _03737_ = \bapg_rd.w_ptr_r [2] ? _03736_ : _03733_;
  assign _03738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [2] : \MSYNC_1r1w.synth.nz.mem[616] [2];
  assign _03739_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [2] : \MSYNC_1r1w.synth.nz.mem[618] [2];
  assign _03740_ = \bapg_rd.w_ptr_r [1] ? _03739_ : _03738_;
  assign _03741_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [2] : \MSYNC_1r1w.synth.nz.mem[620] [2];
  assign _03742_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [2] : \MSYNC_1r1w.synth.nz.mem[622] [2];
  assign _03743_ = \bapg_rd.w_ptr_r [1] ? _03742_ : _03741_;
  assign _03744_ = \bapg_rd.w_ptr_r [2] ? _03743_ : _03740_;
  assign _03745_ = \bapg_rd.w_ptr_r [3] ? _03744_ : _03737_;
  assign _03746_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [2] : \MSYNC_1r1w.synth.nz.mem[624] [2];
  assign _03747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [2] : \MSYNC_1r1w.synth.nz.mem[626] [2];
  assign _03748_ = \bapg_rd.w_ptr_r [1] ? _03747_ : _03746_;
  assign _03749_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [2] : \MSYNC_1r1w.synth.nz.mem[628] [2];
  assign _03750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [2] : \MSYNC_1r1w.synth.nz.mem[630] [2];
  assign _03751_ = \bapg_rd.w_ptr_r [1] ? _03750_ : _03749_;
  assign _03752_ = \bapg_rd.w_ptr_r [2] ? _03751_ : _03748_;
  assign _03753_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [2] : \MSYNC_1r1w.synth.nz.mem[632] [2];
  assign _03754_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [2] : \MSYNC_1r1w.synth.nz.mem[634] [2];
  assign _03755_ = \bapg_rd.w_ptr_r [1] ? _03754_ : _03753_;
  assign _03756_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [2] : \MSYNC_1r1w.synth.nz.mem[636] [2];
  assign _03757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [2] : \MSYNC_1r1w.synth.nz.mem[638] [2];
  assign _03758_ = \bapg_rd.w_ptr_r [1] ? _03757_ : _03756_;
  assign _03759_ = \bapg_rd.w_ptr_r [2] ? _03758_ : _03755_;
  assign _03760_ = \bapg_rd.w_ptr_r [3] ? _03759_ : _03752_;
  assign _03761_ = \bapg_rd.w_ptr_r [4] ? _03760_ : _03745_;
  assign _03762_ = \bapg_rd.w_ptr_r [5] ? _03761_ : _03730_;
  assign _03763_ = \bapg_rd.w_ptr_r [6] ? _03762_ : _03699_;
  assign _03764_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [2] : \MSYNC_1r1w.synth.nz.mem[640] [2];
  assign _03765_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [2] : \MSYNC_1r1w.synth.nz.mem[642] [2];
  assign _03766_ = \bapg_rd.w_ptr_r [1] ? _03765_ : _03764_;
  assign _03767_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [2] : \MSYNC_1r1w.synth.nz.mem[644] [2];
  assign _03768_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [2] : \MSYNC_1r1w.synth.nz.mem[646] [2];
  assign _03769_ = \bapg_rd.w_ptr_r [1] ? _03768_ : _03767_;
  assign _03770_ = \bapg_rd.w_ptr_r [2] ? _03769_ : _03766_;
  assign _03771_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [2] : \MSYNC_1r1w.synth.nz.mem[648] [2];
  assign _03772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [2] : \MSYNC_1r1w.synth.nz.mem[650] [2];
  assign _03773_ = \bapg_rd.w_ptr_r [1] ? _03772_ : _03771_;
  assign _03774_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [2] : \MSYNC_1r1w.synth.nz.mem[652] [2];
  assign _03775_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [2] : \MSYNC_1r1w.synth.nz.mem[654] [2];
  assign _03776_ = \bapg_rd.w_ptr_r [1] ? _03775_ : _03774_;
  assign _03777_ = \bapg_rd.w_ptr_r [2] ? _03776_ : _03773_;
  assign _03778_ = \bapg_rd.w_ptr_r [3] ? _03777_ : _03770_;
  assign _03779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [2] : \MSYNC_1r1w.synth.nz.mem[656] [2];
  assign _03780_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [2] : \MSYNC_1r1w.synth.nz.mem[658] [2];
  assign _03781_ = \bapg_rd.w_ptr_r [1] ? _03780_ : _03779_;
  assign _03782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [2] : \MSYNC_1r1w.synth.nz.mem[660] [2];
  assign _03783_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [2] : \MSYNC_1r1w.synth.nz.mem[662] [2];
  assign _03784_ = \bapg_rd.w_ptr_r [1] ? _03783_ : _03782_;
  assign _03785_ = \bapg_rd.w_ptr_r [2] ? _03784_ : _03781_;
  assign _03786_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [2] : \MSYNC_1r1w.synth.nz.mem[664] [2];
  assign _03787_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [2] : \MSYNC_1r1w.synth.nz.mem[666] [2];
  assign _03788_ = \bapg_rd.w_ptr_r [1] ? _03787_ : _03786_;
  assign _03789_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [2] : \MSYNC_1r1w.synth.nz.mem[668] [2];
  assign _03790_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [2] : \MSYNC_1r1w.synth.nz.mem[670] [2];
  assign _03791_ = \bapg_rd.w_ptr_r [1] ? _03790_ : _03789_;
  assign _03792_ = \bapg_rd.w_ptr_r [2] ? _03791_ : _03788_;
  assign _03793_ = \bapg_rd.w_ptr_r [3] ? _03792_ : _03785_;
  assign _03794_ = \bapg_rd.w_ptr_r [4] ? _03793_ : _03778_;
  assign _03795_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [2] : \MSYNC_1r1w.synth.nz.mem[672] [2];
  assign _03796_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [2] : \MSYNC_1r1w.synth.nz.mem[674] [2];
  assign _03797_ = \bapg_rd.w_ptr_r [1] ? _03796_ : _03795_;
  assign _03798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [2] : \MSYNC_1r1w.synth.nz.mem[676] [2];
  assign _03799_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [2] : \MSYNC_1r1w.synth.nz.mem[678] [2];
  assign _03800_ = \bapg_rd.w_ptr_r [1] ? _03799_ : _03798_;
  assign _03801_ = \bapg_rd.w_ptr_r [2] ? _03800_ : _03797_;
  assign _03802_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [2] : \MSYNC_1r1w.synth.nz.mem[680] [2];
  assign _03803_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [2] : \MSYNC_1r1w.synth.nz.mem[682] [2];
  assign _03804_ = \bapg_rd.w_ptr_r [1] ? _03803_ : _03802_;
  assign _03805_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [2] : \MSYNC_1r1w.synth.nz.mem[684] [2];
  assign _03806_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [2] : \MSYNC_1r1w.synth.nz.mem[686] [2];
  assign _03807_ = \bapg_rd.w_ptr_r [1] ? _03806_ : _03805_;
  assign _03808_ = \bapg_rd.w_ptr_r [2] ? _03807_ : _03804_;
  assign _03809_ = \bapg_rd.w_ptr_r [3] ? _03808_ : _03801_;
  assign _03810_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [2] : \MSYNC_1r1w.synth.nz.mem[688] [2];
  assign _03811_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [2] : \MSYNC_1r1w.synth.nz.mem[690] [2];
  assign _03812_ = \bapg_rd.w_ptr_r [1] ? _03811_ : _03810_;
  assign _03813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [2] : \MSYNC_1r1w.synth.nz.mem[692] [2];
  assign _03814_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [2] : \MSYNC_1r1w.synth.nz.mem[694] [2];
  assign _03815_ = \bapg_rd.w_ptr_r [1] ? _03814_ : _03813_;
  assign _03816_ = \bapg_rd.w_ptr_r [2] ? _03815_ : _03812_;
  assign _03817_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [2] : \MSYNC_1r1w.synth.nz.mem[696] [2];
  assign _03818_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [2] : \MSYNC_1r1w.synth.nz.mem[698] [2];
  assign _03819_ = \bapg_rd.w_ptr_r [1] ? _03818_ : _03817_;
  assign _03820_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [2] : \MSYNC_1r1w.synth.nz.mem[700] [2];
  assign _03821_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [2] : \MSYNC_1r1w.synth.nz.mem[702] [2];
  assign _03822_ = \bapg_rd.w_ptr_r [1] ? _03821_ : _03820_;
  assign _03823_ = \bapg_rd.w_ptr_r [2] ? _03822_ : _03819_;
  assign _03824_ = \bapg_rd.w_ptr_r [3] ? _03823_ : _03816_;
  assign _03825_ = \bapg_rd.w_ptr_r [4] ? _03824_ : _03809_;
  assign _03826_ = \bapg_rd.w_ptr_r [5] ? _03825_ : _03794_;
  assign _03827_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [2] : \MSYNC_1r1w.synth.nz.mem[704] [2];
  assign _03828_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [2] : \MSYNC_1r1w.synth.nz.mem[706] [2];
  assign _03829_ = \bapg_rd.w_ptr_r [1] ? _03828_ : _03827_;
  assign _03830_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [2] : \MSYNC_1r1w.synth.nz.mem[708] [2];
  assign _03831_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [2] : \MSYNC_1r1w.synth.nz.mem[710] [2];
  assign _03832_ = \bapg_rd.w_ptr_r [1] ? _03831_ : _03830_;
  assign _03833_ = \bapg_rd.w_ptr_r [2] ? _03832_ : _03829_;
  assign _03834_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [2] : \MSYNC_1r1w.synth.nz.mem[712] [2];
  assign _03835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [2] : \MSYNC_1r1w.synth.nz.mem[714] [2];
  assign _03836_ = \bapg_rd.w_ptr_r [1] ? _03835_ : _03834_;
  assign _03837_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [2] : \MSYNC_1r1w.synth.nz.mem[716] [2];
  assign _03838_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [2] : \MSYNC_1r1w.synth.nz.mem[718] [2];
  assign _03839_ = \bapg_rd.w_ptr_r [1] ? _03838_ : _03837_;
  assign _03840_ = \bapg_rd.w_ptr_r [2] ? _03839_ : _03836_;
  assign _03841_ = \bapg_rd.w_ptr_r [3] ? _03840_ : _03833_;
  assign _03842_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [2] : \MSYNC_1r1w.synth.nz.mem[720] [2];
  assign _03843_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [2] : \MSYNC_1r1w.synth.nz.mem[722] [2];
  assign _03844_ = \bapg_rd.w_ptr_r [1] ? _03843_ : _03842_;
  assign _03845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [2] : \MSYNC_1r1w.synth.nz.mem[724] [2];
  assign _03846_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [2] : \MSYNC_1r1w.synth.nz.mem[726] [2];
  assign _03847_ = \bapg_rd.w_ptr_r [1] ? _03846_ : _03845_;
  assign _03848_ = \bapg_rd.w_ptr_r [2] ? _03847_ : _03844_;
  assign _03849_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [2] : \MSYNC_1r1w.synth.nz.mem[728] [2];
  assign _03850_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [2] : \MSYNC_1r1w.synth.nz.mem[730] [2];
  assign _03851_ = \bapg_rd.w_ptr_r [1] ? _03850_ : _03849_;
  assign _03852_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [2] : \MSYNC_1r1w.synth.nz.mem[732] [2];
  assign _03853_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [2] : \MSYNC_1r1w.synth.nz.mem[734] [2];
  assign _03854_ = \bapg_rd.w_ptr_r [1] ? _03853_ : _03852_;
  assign _03855_ = \bapg_rd.w_ptr_r [2] ? _03854_ : _03851_;
  assign _03856_ = \bapg_rd.w_ptr_r [3] ? _03855_ : _03848_;
  assign _03857_ = \bapg_rd.w_ptr_r [4] ? _03856_ : _03841_;
  assign _03858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [2] : \MSYNC_1r1w.synth.nz.mem[736] [2];
  assign _03859_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [2] : \MSYNC_1r1w.synth.nz.mem[738] [2];
  assign _03860_ = \bapg_rd.w_ptr_r [1] ? _03859_ : _03858_;
  assign _03861_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [2] : \MSYNC_1r1w.synth.nz.mem[740] [2];
  assign _03862_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [2] : \MSYNC_1r1w.synth.nz.mem[742] [2];
  assign _03863_ = \bapg_rd.w_ptr_r [1] ? _03862_ : _03861_;
  assign _03864_ = \bapg_rd.w_ptr_r [2] ? _03863_ : _03860_;
  assign _03865_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [2] : \MSYNC_1r1w.synth.nz.mem[744] [2];
  assign _03866_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [2] : \MSYNC_1r1w.synth.nz.mem[746] [2];
  assign _03867_ = \bapg_rd.w_ptr_r [1] ? _03866_ : _03865_;
  assign _03868_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [2] : \MSYNC_1r1w.synth.nz.mem[748] [2];
  assign _03869_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [2] : \MSYNC_1r1w.synth.nz.mem[750] [2];
  assign _03870_ = \bapg_rd.w_ptr_r [1] ? _03869_ : _03868_;
  assign _03871_ = \bapg_rd.w_ptr_r [2] ? _03870_ : _03867_;
  assign _03872_ = \bapg_rd.w_ptr_r [3] ? _03871_ : _03864_;
  assign _03873_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [2] : \MSYNC_1r1w.synth.nz.mem[752] [2];
  assign _03874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [2] : \MSYNC_1r1w.synth.nz.mem[754] [2];
  assign _03875_ = \bapg_rd.w_ptr_r [1] ? _03874_ : _03873_;
  assign _03876_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [2] : \MSYNC_1r1w.synth.nz.mem[756] [2];
  assign _03877_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [2] : \MSYNC_1r1w.synth.nz.mem[758] [2];
  assign _03878_ = \bapg_rd.w_ptr_r [1] ? _03877_ : _03876_;
  assign _03879_ = \bapg_rd.w_ptr_r [2] ? _03878_ : _03875_;
  assign _03880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [2] : \MSYNC_1r1w.synth.nz.mem[760] [2];
  assign _03881_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [2] : \MSYNC_1r1w.synth.nz.mem[762] [2];
  assign _03882_ = \bapg_rd.w_ptr_r [1] ? _03881_ : _03880_;
  assign _03883_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [2] : \MSYNC_1r1w.synth.nz.mem[764] [2];
  assign _03884_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [2] : \MSYNC_1r1w.synth.nz.mem[766] [2];
  assign _03885_ = \bapg_rd.w_ptr_r [1] ? _03884_ : _03883_;
  assign _03886_ = \bapg_rd.w_ptr_r [2] ? _03885_ : _03882_;
  assign _03887_ = \bapg_rd.w_ptr_r [3] ? _03886_ : _03879_;
  assign _03888_ = \bapg_rd.w_ptr_r [4] ? _03887_ : _03872_;
  assign _03889_ = \bapg_rd.w_ptr_r [5] ? _03888_ : _03857_;
  assign _03890_ = \bapg_rd.w_ptr_r [6] ? _03889_ : _03826_;
  assign _03891_ = \bapg_rd.w_ptr_r [7] ? _03890_ : _03763_;
  assign _03892_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [2] : \MSYNC_1r1w.synth.nz.mem[768] [2];
  assign _03893_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [2] : \MSYNC_1r1w.synth.nz.mem[770] [2];
  assign _03894_ = \bapg_rd.w_ptr_r [1] ? _03893_ : _03892_;
  assign _03895_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [2] : \MSYNC_1r1w.synth.nz.mem[772] [2];
  assign _03896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [2] : \MSYNC_1r1w.synth.nz.mem[774] [2];
  assign _03897_ = \bapg_rd.w_ptr_r [1] ? _03896_ : _03895_;
  assign _03898_ = \bapg_rd.w_ptr_r [2] ? _03897_ : _03894_;
  assign _03899_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [2] : \MSYNC_1r1w.synth.nz.mem[776] [2];
  assign _03900_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [2] : \MSYNC_1r1w.synth.nz.mem[778] [2];
  assign _03901_ = \bapg_rd.w_ptr_r [1] ? _03900_ : _03899_;
  assign _03902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [2] : \MSYNC_1r1w.synth.nz.mem[780] [2];
  assign _03903_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [2] : \MSYNC_1r1w.synth.nz.mem[782] [2];
  assign _03904_ = \bapg_rd.w_ptr_r [1] ? _03903_ : _03902_;
  assign _03905_ = \bapg_rd.w_ptr_r [2] ? _03904_ : _03901_;
  assign _03906_ = \bapg_rd.w_ptr_r [3] ? _03905_ : _03898_;
  assign _03907_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [2] : \MSYNC_1r1w.synth.nz.mem[784] [2];
  assign _03908_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [2] : \MSYNC_1r1w.synth.nz.mem[786] [2];
  assign _03909_ = \bapg_rd.w_ptr_r [1] ? _03908_ : _03907_;
  assign _03910_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [2] : \MSYNC_1r1w.synth.nz.mem[788] [2];
  assign _03911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [2] : \MSYNC_1r1w.synth.nz.mem[790] [2];
  assign _03912_ = \bapg_rd.w_ptr_r [1] ? _03911_ : _03910_;
  assign _03913_ = \bapg_rd.w_ptr_r [2] ? _03912_ : _03909_;
  assign _03914_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [2] : \MSYNC_1r1w.synth.nz.mem[792] [2];
  assign _03915_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [2] : \MSYNC_1r1w.synth.nz.mem[794] [2];
  assign _03916_ = \bapg_rd.w_ptr_r [1] ? _03915_ : _03914_;
  assign _03917_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [2] : \MSYNC_1r1w.synth.nz.mem[796] [2];
  assign _03918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [2] : \MSYNC_1r1w.synth.nz.mem[798] [2];
  assign _03919_ = \bapg_rd.w_ptr_r [1] ? _03918_ : _03917_;
  assign _03920_ = \bapg_rd.w_ptr_r [2] ? _03919_ : _03916_;
  assign _03921_ = \bapg_rd.w_ptr_r [3] ? _03920_ : _03913_;
  assign _03922_ = \bapg_rd.w_ptr_r [4] ? _03921_ : _03906_;
  assign _03923_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [2] : \MSYNC_1r1w.synth.nz.mem[800] [2];
  assign _03924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [2] : \MSYNC_1r1w.synth.nz.mem[802] [2];
  assign _03925_ = \bapg_rd.w_ptr_r [1] ? _03924_ : _03923_;
  assign _03926_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [2] : \MSYNC_1r1w.synth.nz.mem[804] [2];
  assign _03927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [2] : \MSYNC_1r1w.synth.nz.mem[806] [2];
  assign _03928_ = \bapg_rd.w_ptr_r [1] ? _03927_ : _03926_;
  assign _03929_ = \bapg_rd.w_ptr_r [2] ? _03928_ : _03925_;
  assign _03930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [2] : \MSYNC_1r1w.synth.nz.mem[808] [2];
  assign _03931_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [2] : \MSYNC_1r1w.synth.nz.mem[810] [2];
  assign _03932_ = \bapg_rd.w_ptr_r [1] ? _03931_ : _03930_;
  assign _03933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [2] : \MSYNC_1r1w.synth.nz.mem[812] [2];
  assign _03934_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [2] : \MSYNC_1r1w.synth.nz.mem[814] [2];
  assign _03935_ = \bapg_rd.w_ptr_r [1] ? _03934_ : _03933_;
  assign _03936_ = \bapg_rd.w_ptr_r [2] ? _03935_ : _03932_;
  assign _03937_ = \bapg_rd.w_ptr_r [3] ? _03936_ : _03929_;
  assign _03938_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [2] : \MSYNC_1r1w.synth.nz.mem[816] [2];
  assign _03939_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [2] : \MSYNC_1r1w.synth.nz.mem[818] [2];
  assign _03940_ = \bapg_rd.w_ptr_r [1] ? _03939_ : _03938_;
  assign _03941_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [2] : \MSYNC_1r1w.synth.nz.mem[820] [2];
  assign _03942_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [2] : \MSYNC_1r1w.synth.nz.mem[822] [2];
  assign _03943_ = \bapg_rd.w_ptr_r [1] ? _03942_ : _03941_;
  assign _03944_ = \bapg_rd.w_ptr_r [2] ? _03943_ : _03940_;
  assign _03945_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [2] : \MSYNC_1r1w.synth.nz.mem[824] [2];
  assign _03946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [2] : \MSYNC_1r1w.synth.nz.mem[826] [2];
  assign _03947_ = \bapg_rd.w_ptr_r [1] ? _03946_ : _03945_;
  assign _03948_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [2] : \MSYNC_1r1w.synth.nz.mem[828] [2];
  assign _03949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [2] : \MSYNC_1r1w.synth.nz.mem[830] [2];
  assign _03950_ = \bapg_rd.w_ptr_r [1] ? _03949_ : _03948_;
  assign _03951_ = \bapg_rd.w_ptr_r [2] ? _03950_ : _03947_;
  assign _03952_ = \bapg_rd.w_ptr_r [3] ? _03951_ : _03944_;
  assign _03953_ = \bapg_rd.w_ptr_r [4] ? _03952_ : _03937_;
  assign _03954_ = \bapg_rd.w_ptr_r [5] ? _03953_ : _03922_;
  assign _03955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [2] : \MSYNC_1r1w.synth.nz.mem[832] [2];
  assign _03956_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [2] : \MSYNC_1r1w.synth.nz.mem[834] [2];
  assign _03957_ = \bapg_rd.w_ptr_r [1] ? _03956_ : _03955_;
  assign _03958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [2] : \MSYNC_1r1w.synth.nz.mem[836] [2];
  assign _03959_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [2] : \MSYNC_1r1w.synth.nz.mem[838] [2];
  assign _03960_ = \bapg_rd.w_ptr_r [1] ? _03959_ : _03958_;
  assign _03961_ = \bapg_rd.w_ptr_r [2] ? _03960_ : _03957_;
  assign _03962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [2] : \MSYNC_1r1w.synth.nz.mem[840] [2];
  assign _03963_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [2] : \MSYNC_1r1w.synth.nz.mem[842] [2];
  assign _03964_ = \bapg_rd.w_ptr_r [1] ? _03963_ : _03962_;
  assign _03965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [2] : \MSYNC_1r1w.synth.nz.mem[844] [2];
  assign _03966_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [2] : \MSYNC_1r1w.synth.nz.mem[846] [2];
  assign _03967_ = \bapg_rd.w_ptr_r [1] ? _03966_ : _03965_;
  assign _03968_ = \bapg_rd.w_ptr_r [2] ? _03967_ : _03964_;
  assign _03969_ = \bapg_rd.w_ptr_r [3] ? _03968_ : _03961_;
  assign _03970_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [2] : \MSYNC_1r1w.synth.nz.mem[848] [2];
  assign _03971_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [2] : \MSYNC_1r1w.synth.nz.mem[850] [2];
  assign _03972_ = \bapg_rd.w_ptr_r [1] ? _03971_ : _03970_;
  assign _03973_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [2] : \MSYNC_1r1w.synth.nz.mem[852] [2];
  assign _03974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [2] : \MSYNC_1r1w.synth.nz.mem[854] [2];
  assign _03975_ = \bapg_rd.w_ptr_r [1] ? _03974_ : _03973_;
  assign _03976_ = \bapg_rd.w_ptr_r [2] ? _03975_ : _03972_;
  assign _03977_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [2] : \MSYNC_1r1w.synth.nz.mem[856] [2];
  assign _03978_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [2] : \MSYNC_1r1w.synth.nz.mem[858] [2];
  assign _03979_ = \bapg_rd.w_ptr_r [1] ? _03978_ : _03977_;
  assign _03980_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [2] : \MSYNC_1r1w.synth.nz.mem[860] [2];
  assign _03981_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [2] : \MSYNC_1r1w.synth.nz.mem[862] [2];
  assign _03982_ = \bapg_rd.w_ptr_r [1] ? _03981_ : _03980_;
  assign _03983_ = \bapg_rd.w_ptr_r [2] ? _03982_ : _03979_;
  assign _03984_ = \bapg_rd.w_ptr_r [3] ? _03983_ : _03976_;
  assign _03985_ = \bapg_rd.w_ptr_r [4] ? _03984_ : _03969_;
  assign _03986_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [2] : \MSYNC_1r1w.synth.nz.mem[864] [2];
  assign _03987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [2] : \MSYNC_1r1w.synth.nz.mem[866] [2];
  assign _03988_ = \bapg_rd.w_ptr_r [1] ? _03987_ : _03986_;
  assign _03989_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [2] : \MSYNC_1r1w.synth.nz.mem[868] [2];
  assign _03990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [2] : \MSYNC_1r1w.synth.nz.mem[870] [2];
  assign _03991_ = \bapg_rd.w_ptr_r [1] ? _03990_ : _03989_;
  assign _03992_ = \bapg_rd.w_ptr_r [2] ? _03991_ : _03988_;
  assign _03993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [2] : \MSYNC_1r1w.synth.nz.mem[872] [2];
  assign _03994_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [2] : \MSYNC_1r1w.synth.nz.mem[874] [2];
  assign _03995_ = \bapg_rd.w_ptr_r [1] ? _03994_ : _03993_;
  assign _03996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [2] : \MSYNC_1r1w.synth.nz.mem[876] [2];
  assign _03997_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [2] : \MSYNC_1r1w.synth.nz.mem[878] [2];
  assign _03998_ = \bapg_rd.w_ptr_r [1] ? _03997_ : _03996_;
  assign _03999_ = \bapg_rd.w_ptr_r [2] ? _03998_ : _03995_;
  assign _04000_ = \bapg_rd.w_ptr_r [3] ? _03999_ : _03992_;
  assign _04001_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [2] : \MSYNC_1r1w.synth.nz.mem[880] [2];
  assign _04002_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [2] : \MSYNC_1r1w.synth.nz.mem[882] [2];
  assign _04003_ = \bapg_rd.w_ptr_r [1] ? _04002_ : _04001_;
  assign _04004_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [2] : \MSYNC_1r1w.synth.nz.mem[884] [2];
  assign _04005_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [2] : \MSYNC_1r1w.synth.nz.mem[886] [2];
  assign _04006_ = \bapg_rd.w_ptr_r [1] ? _04005_ : _04004_;
  assign _04007_ = \bapg_rd.w_ptr_r [2] ? _04006_ : _04003_;
  assign _04008_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [2] : \MSYNC_1r1w.synth.nz.mem[888] [2];
  assign _04009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [2] : \MSYNC_1r1w.synth.nz.mem[890] [2];
  assign _04010_ = \bapg_rd.w_ptr_r [1] ? _04009_ : _04008_;
  assign _04011_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [2] : \MSYNC_1r1w.synth.nz.mem[892] [2];
  assign _04012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [2] : \MSYNC_1r1w.synth.nz.mem[894] [2];
  assign _04013_ = \bapg_rd.w_ptr_r [1] ? _04012_ : _04011_;
  assign _04014_ = \bapg_rd.w_ptr_r [2] ? _04013_ : _04010_;
  assign _04015_ = \bapg_rd.w_ptr_r [3] ? _04014_ : _04007_;
  assign _04016_ = \bapg_rd.w_ptr_r [4] ? _04015_ : _04000_;
  assign _04017_ = \bapg_rd.w_ptr_r [5] ? _04016_ : _03985_;
  assign _04018_ = \bapg_rd.w_ptr_r [6] ? _04017_ : _03954_;
  assign _04019_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [2] : \MSYNC_1r1w.synth.nz.mem[896] [2];
  assign _04020_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [2] : \MSYNC_1r1w.synth.nz.mem[898] [2];
  assign _04021_ = \bapg_rd.w_ptr_r [1] ? _04020_ : _04019_;
  assign _04022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [2] : \MSYNC_1r1w.synth.nz.mem[900] [2];
  assign _04023_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [2] : \MSYNC_1r1w.synth.nz.mem[902] [2];
  assign _04024_ = \bapg_rd.w_ptr_r [1] ? _04023_ : _04022_;
  assign _04025_ = \bapg_rd.w_ptr_r [2] ? _04024_ : _04021_;
  assign _04026_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [2] : \MSYNC_1r1w.synth.nz.mem[904] [2];
  assign _04027_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [2] : \MSYNC_1r1w.synth.nz.mem[906] [2];
  assign _04028_ = \bapg_rd.w_ptr_r [1] ? _04027_ : _04026_;
  assign _04029_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [2] : \MSYNC_1r1w.synth.nz.mem[908] [2];
  assign _04030_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [2] : \MSYNC_1r1w.synth.nz.mem[910] [2];
  assign _04031_ = \bapg_rd.w_ptr_r [1] ? _04030_ : _04029_;
  assign _04032_ = \bapg_rd.w_ptr_r [2] ? _04031_ : _04028_;
  assign _04033_ = \bapg_rd.w_ptr_r [3] ? _04032_ : _04025_;
  assign _04034_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [2] : \MSYNC_1r1w.synth.nz.mem[912] [2];
  assign _04035_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [2] : \MSYNC_1r1w.synth.nz.mem[914] [2];
  assign _04036_ = \bapg_rd.w_ptr_r [1] ? _04035_ : _04034_;
  assign _04037_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [2] : \MSYNC_1r1w.synth.nz.mem[916] [2];
  assign _04038_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [2] : \MSYNC_1r1w.synth.nz.mem[918] [2];
  assign _04039_ = \bapg_rd.w_ptr_r [1] ? _04038_ : _04037_;
  assign _04040_ = \bapg_rd.w_ptr_r [2] ? _04039_ : _04036_;
  assign _04041_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [2] : \MSYNC_1r1w.synth.nz.mem[920] [2];
  assign _04042_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [2] : \MSYNC_1r1w.synth.nz.mem[922] [2];
  assign _04043_ = \bapg_rd.w_ptr_r [1] ? _04042_ : _04041_;
  assign _04044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [2] : \MSYNC_1r1w.synth.nz.mem[924] [2];
  assign _04045_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [2] : \MSYNC_1r1w.synth.nz.mem[926] [2];
  assign _04046_ = \bapg_rd.w_ptr_r [1] ? _04045_ : _04044_;
  assign _04047_ = \bapg_rd.w_ptr_r [2] ? _04046_ : _04043_;
  assign _04048_ = \bapg_rd.w_ptr_r [3] ? _04047_ : _04040_;
  assign _04049_ = \bapg_rd.w_ptr_r [4] ? _04048_ : _04033_;
  assign _04050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [2] : \MSYNC_1r1w.synth.nz.mem[928] [2];
  assign _04051_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [2] : \MSYNC_1r1w.synth.nz.mem[930] [2];
  assign _04052_ = \bapg_rd.w_ptr_r [1] ? _04051_ : _04050_;
  assign _04053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [2] : \MSYNC_1r1w.synth.nz.mem[932] [2];
  assign _04054_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [2] : \MSYNC_1r1w.synth.nz.mem[934] [2];
  assign _04055_ = \bapg_rd.w_ptr_r [1] ? _04054_ : _04053_;
  assign _04056_ = \bapg_rd.w_ptr_r [2] ? _04055_ : _04052_;
  assign _04057_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [2] : \MSYNC_1r1w.synth.nz.mem[936] [2];
  assign _04058_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [2] : \MSYNC_1r1w.synth.nz.mem[938] [2];
  assign _04059_ = \bapg_rd.w_ptr_r [1] ? _04058_ : _04057_;
  assign _04060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [2] : \MSYNC_1r1w.synth.nz.mem[940] [2];
  assign _04061_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [2] : \MSYNC_1r1w.synth.nz.mem[942] [2];
  assign _04062_ = \bapg_rd.w_ptr_r [1] ? _04061_ : _04060_;
  assign _04063_ = \bapg_rd.w_ptr_r [2] ? _04062_ : _04059_;
  assign _04064_ = \bapg_rd.w_ptr_r [3] ? _04063_ : _04056_;
  assign _04065_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [2] : \MSYNC_1r1w.synth.nz.mem[944] [2];
  assign _04066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [2] : \MSYNC_1r1w.synth.nz.mem[946] [2];
  assign _04067_ = \bapg_rd.w_ptr_r [1] ? _04066_ : _04065_;
  assign _04068_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [2] : \MSYNC_1r1w.synth.nz.mem[948] [2];
  assign _04069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [2] : \MSYNC_1r1w.synth.nz.mem[950] [2];
  assign _04070_ = \bapg_rd.w_ptr_r [1] ? _04069_ : _04068_;
  assign _04071_ = \bapg_rd.w_ptr_r [2] ? _04070_ : _04067_;
  assign _04072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [2] : \MSYNC_1r1w.synth.nz.mem[952] [2];
  assign _04073_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [2] : \MSYNC_1r1w.synth.nz.mem[954] [2];
  assign _04074_ = \bapg_rd.w_ptr_r [1] ? _04073_ : _04072_;
  assign _04075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [2] : \MSYNC_1r1w.synth.nz.mem[956] [2];
  assign _04076_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [2] : \MSYNC_1r1w.synth.nz.mem[958] [2];
  assign _04077_ = \bapg_rd.w_ptr_r [1] ? _04076_ : _04075_;
  assign _04078_ = \bapg_rd.w_ptr_r [2] ? _04077_ : _04074_;
  assign _04079_ = \bapg_rd.w_ptr_r [3] ? _04078_ : _04071_;
  assign _04080_ = \bapg_rd.w_ptr_r [4] ? _04079_ : _04064_;
  assign _04081_ = \bapg_rd.w_ptr_r [5] ? _04080_ : _04049_;
  assign _04082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [2] : \MSYNC_1r1w.synth.nz.mem[960] [2];
  assign _04083_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [2] : \MSYNC_1r1w.synth.nz.mem[962] [2];
  assign _04084_ = \bapg_rd.w_ptr_r [1] ? _04083_ : _04082_;
  assign _04085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [2] : \MSYNC_1r1w.synth.nz.mem[964] [2];
  assign _04086_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [2] : \MSYNC_1r1w.synth.nz.mem[966] [2];
  assign _04087_ = \bapg_rd.w_ptr_r [1] ? _04086_ : _04085_;
  assign _04088_ = \bapg_rd.w_ptr_r [2] ? _04087_ : _04084_;
  assign _04089_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [2] : \MSYNC_1r1w.synth.nz.mem[968] [2];
  assign _04090_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [2] : \MSYNC_1r1w.synth.nz.mem[970] [2];
  assign _04091_ = \bapg_rd.w_ptr_r [1] ? _04090_ : _04089_;
  assign _04092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [2] : \MSYNC_1r1w.synth.nz.mem[972] [2];
  assign _04093_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [2] : \MSYNC_1r1w.synth.nz.mem[974] [2];
  assign _04094_ = \bapg_rd.w_ptr_r [1] ? _04093_ : _04092_;
  assign _04095_ = \bapg_rd.w_ptr_r [2] ? _04094_ : _04091_;
  assign _04096_ = \bapg_rd.w_ptr_r [3] ? _04095_ : _04088_;
  assign _04097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [2] : \MSYNC_1r1w.synth.nz.mem[976] [2];
  assign _04098_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [2] : \MSYNC_1r1w.synth.nz.mem[978] [2];
  assign _04099_ = \bapg_rd.w_ptr_r [1] ? _04098_ : _04097_;
  assign _04100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [2] : \MSYNC_1r1w.synth.nz.mem[980] [2];
  assign _04101_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [2] : \MSYNC_1r1w.synth.nz.mem[982] [2];
  assign _04102_ = \bapg_rd.w_ptr_r [1] ? _04101_ : _04100_;
  assign _04103_ = \bapg_rd.w_ptr_r [2] ? _04102_ : _04099_;
  assign _04104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [2] : \MSYNC_1r1w.synth.nz.mem[984] [2];
  assign _04105_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [2] : \MSYNC_1r1w.synth.nz.mem[986] [2];
  assign _04106_ = \bapg_rd.w_ptr_r [1] ? _04105_ : _04104_;
  assign _04107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [2] : \MSYNC_1r1w.synth.nz.mem[988] [2];
  assign _04108_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [2] : \MSYNC_1r1w.synth.nz.mem[990] [2];
  assign _04109_ = \bapg_rd.w_ptr_r [1] ? _04108_ : _04107_;
  assign _04110_ = \bapg_rd.w_ptr_r [2] ? _04109_ : _04106_;
  assign _04111_ = \bapg_rd.w_ptr_r [3] ? _04110_ : _04103_;
  assign _04112_ = \bapg_rd.w_ptr_r [4] ? _04111_ : _04096_;
  assign _04113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [2] : \MSYNC_1r1w.synth.nz.mem[992] [2];
  assign _04114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [2] : \MSYNC_1r1w.synth.nz.mem[994] [2];
  assign _04115_ = \bapg_rd.w_ptr_r [1] ? _04114_ : _04113_;
  assign _04116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [2] : \MSYNC_1r1w.synth.nz.mem[996] [2];
  assign _04117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [2] : \MSYNC_1r1w.synth.nz.mem[998] [2];
  assign _04118_ = \bapg_rd.w_ptr_r [1] ? _04117_ : _04116_;
  assign _04119_ = \bapg_rd.w_ptr_r [2] ? _04118_ : _04115_;
  assign _04120_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [2] : \MSYNC_1r1w.synth.nz.mem[1000] [2];
  assign _04121_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [2] : \MSYNC_1r1w.synth.nz.mem[1002] [2];
  assign _04122_ = \bapg_rd.w_ptr_r [1] ? _04121_ : _04120_;
  assign _04123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [2] : \MSYNC_1r1w.synth.nz.mem[1004] [2];
  assign _04124_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [2] : \MSYNC_1r1w.synth.nz.mem[1006] [2];
  assign _04125_ = \bapg_rd.w_ptr_r [1] ? _04124_ : _04123_;
  assign _04126_ = \bapg_rd.w_ptr_r [2] ? _04125_ : _04122_;
  assign _04127_ = \bapg_rd.w_ptr_r [3] ? _04126_ : _04119_;
  assign _04128_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [2] : \MSYNC_1r1w.synth.nz.mem[1008] [2];
  assign _04129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [2] : \MSYNC_1r1w.synth.nz.mem[1010] [2];
  assign _04130_ = \bapg_rd.w_ptr_r [1] ? _04129_ : _04128_;
  assign _04131_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [2] : \MSYNC_1r1w.synth.nz.mem[1012] [2];
  assign _04132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [2] : \MSYNC_1r1w.synth.nz.mem[1014] [2];
  assign _04133_ = \bapg_rd.w_ptr_r [1] ? _04132_ : _04131_;
  assign _04134_ = \bapg_rd.w_ptr_r [2] ? _04133_ : _04130_;
  assign _04135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [2] : \MSYNC_1r1w.synth.nz.mem[1016] [2];
  assign _04136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [2] : \MSYNC_1r1w.synth.nz.mem[1018] [2];
  assign _04137_ = \bapg_rd.w_ptr_r [1] ? _04136_ : _04135_;
  assign _04138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [2] : \MSYNC_1r1w.synth.nz.mem[1020] [2];
  assign _04139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [2] : \MSYNC_1r1w.synth.nz.mem[1022] [2];
  assign _04140_ = \bapg_rd.w_ptr_r [1] ? _04139_ : _04138_;
  assign _04141_ = \bapg_rd.w_ptr_r [2] ? _04140_ : _04137_;
  assign _04142_ = \bapg_rd.w_ptr_r [3] ? _04141_ : _04134_;
  assign _04143_ = \bapg_rd.w_ptr_r [4] ? _04142_ : _04127_;
  assign _04144_ = \bapg_rd.w_ptr_r [5] ? _04143_ : _04112_;
  assign _04145_ = \bapg_rd.w_ptr_r [6] ? _04144_ : _04081_;
  assign _04146_ = \bapg_rd.w_ptr_r [7] ? _04145_ : _04018_;
  assign _04147_ = \bapg_rd.w_ptr_r [8] ? _04146_ : _03891_;
  assign r_data_o[2] = \bapg_rd.w_ptr_r [9] ? _04147_ : _03636_;
  assign _04148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [3] : \MSYNC_1r1w.synth.nz.mem[0] [3];
  assign _04149_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [3] : \MSYNC_1r1w.synth.nz.mem[2] [3];
  assign _04150_ = \bapg_rd.w_ptr_r [1] ? _04149_ : _04148_;
  assign _04151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [3] : \MSYNC_1r1w.synth.nz.mem[4] [3];
  assign _04152_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [3] : \MSYNC_1r1w.synth.nz.mem[6] [3];
  assign _04153_ = \bapg_rd.w_ptr_r [1] ? _04152_ : _04151_;
  assign _04154_ = \bapg_rd.w_ptr_r [2] ? _04153_ : _04150_;
  assign _04155_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [3] : \MSYNC_1r1w.synth.nz.mem[8] [3];
  assign _04156_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [3] : \MSYNC_1r1w.synth.nz.mem[10] [3];
  assign _04157_ = \bapg_rd.w_ptr_r [1] ? _04156_ : _04155_;
  assign _04158_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [3] : \MSYNC_1r1w.synth.nz.mem[12] [3];
  assign _04159_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [3] : \MSYNC_1r1w.synth.nz.mem[14] [3];
  assign _04160_ = \bapg_rd.w_ptr_r [1] ? _04159_ : _04158_;
  assign _04161_ = \bapg_rd.w_ptr_r [2] ? _04160_ : _04157_;
  assign _04162_ = \bapg_rd.w_ptr_r [3] ? _04161_ : _04154_;
  assign _04163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [3] : \MSYNC_1r1w.synth.nz.mem[16] [3];
  assign _04164_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [3] : \MSYNC_1r1w.synth.nz.mem[18] [3];
  assign _04165_ = \bapg_rd.w_ptr_r [1] ? _04164_ : _04163_;
  assign _04166_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [3] : \MSYNC_1r1w.synth.nz.mem[20] [3];
  assign _04167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [3] : \MSYNC_1r1w.synth.nz.mem[22] [3];
  assign _04168_ = \bapg_rd.w_ptr_r [1] ? _04167_ : _04166_;
  assign _04169_ = \bapg_rd.w_ptr_r [2] ? _04168_ : _04165_;
  assign _04170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [3] : \MSYNC_1r1w.synth.nz.mem[24] [3];
  assign _04171_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [3] : \MSYNC_1r1w.synth.nz.mem[26] [3];
  assign _04172_ = \bapg_rd.w_ptr_r [1] ? _04171_ : _04170_;
  assign _04173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [3] : \MSYNC_1r1w.synth.nz.mem[28] [3];
  assign _04174_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [3] : \MSYNC_1r1w.synth.nz.mem[30] [3];
  assign _04175_ = \bapg_rd.w_ptr_r [1] ? _04174_ : _04173_;
  assign _04176_ = \bapg_rd.w_ptr_r [2] ? _04175_ : _04172_;
  assign _04177_ = \bapg_rd.w_ptr_r [3] ? _04176_ : _04169_;
  assign _04178_ = \bapg_rd.w_ptr_r [4] ? _04177_ : _04162_;
  assign _04179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [3] : \MSYNC_1r1w.synth.nz.mem[32] [3];
  assign _04180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [3] : \MSYNC_1r1w.synth.nz.mem[34] [3];
  assign _04181_ = \bapg_rd.w_ptr_r [1] ? _04180_ : _04179_;
  assign _04182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [3] : \MSYNC_1r1w.synth.nz.mem[36] [3];
  assign _04183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [3] : \MSYNC_1r1w.synth.nz.mem[38] [3];
  assign _04184_ = \bapg_rd.w_ptr_r [1] ? _04183_ : _04182_;
  assign _04185_ = \bapg_rd.w_ptr_r [2] ? _04184_ : _04181_;
  assign _04186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [3] : \MSYNC_1r1w.synth.nz.mem[40] [3];
  assign _04187_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [3] : \MSYNC_1r1w.synth.nz.mem[42] [3];
  assign _04188_ = \bapg_rd.w_ptr_r [1] ? _04187_ : _04186_;
  assign _04189_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [3] : \MSYNC_1r1w.synth.nz.mem[44] [3];
  assign _04190_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [3] : \MSYNC_1r1w.synth.nz.mem[46] [3];
  assign _04191_ = \bapg_rd.w_ptr_r [1] ? _04190_ : _04189_;
  assign _04192_ = \bapg_rd.w_ptr_r [2] ? _04191_ : _04188_;
  assign _04193_ = \bapg_rd.w_ptr_r [3] ? _04192_ : _04185_;
  assign _04194_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [3] : \MSYNC_1r1w.synth.nz.mem[48] [3];
  assign _04195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [3] : \MSYNC_1r1w.synth.nz.mem[50] [3];
  assign _04196_ = \bapg_rd.w_ptr_r [1] ? _04195_ : _04194_;
  assign _04197_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [3] : \MSYNC_1r1w.synth.nz.mem[52] [3];
  assign _04198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [3] : \MSYNC_1r1w.synth.nz.mem[54] [3];
  assign _04199_ = \bapg_rd.w_ptr_r [1] ? _04198_ : _04197_;
  assign _04200_ = \bapg_rd.w_ptr_r [2] ? _04199_ : _04196_;
  assign _04201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [3] : \MSYNC_1r1w.synth.nz.mem[56] [3];
  assign _04202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [3] : \MSYNC_1r1w.synth.nz.mem[58] [3];
  assign _04203_ = \bapg_rd.w_ptr_r [1] ? _04202_ : _04201_;
  assign _04204_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [3] : \MSYNC_1r1w.synth.nz.mem[60] [3];
  assign _04205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [3] : \MSYNC_1r1w.synth.nz.mem[62] [3];
  assign _04206_ = \bapg_rd.w_ptr_r [1] ? _04205_ : _04204_;
  assign _04207_ = \bapg_rd.w_ptr_r [2] ? _04206_ : _04203_;
  assign _04208_ = \bapg_rd.w_ptr_r [3] ? _04207_ : _04200_;
  assign _04209_ = \bapg_rd.w_ptr_r [4] ? _04208_ : _04193_;
  assign _04210_ = \bapg_rd.w_ptr_r [5] ? _04209_ : _04178_;
  assign _04211_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [3] : \MSYNC_1r1w.synth.nz.mem[64] [3];
  assign _04212_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [3] : \MSYNC_1r1w.synth.nz.mem[66] [3];
  assign _04213_ = \bapg_rd.w_ptr_r [1] ? _04212_ : _04211_;
  assign _04214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [3] : \MSYNC_1r1w.synth.nz.mem[68] [3];
  assign _04215_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [3] : \MSYNC_1r1w.synth.nz.mem[70] [3];
  assign _04216_ = \bapg_rd.w_ptr_r [1] ? _04215_ : _04214_;
  assign _04217_ = \bapg_rd.w_ptr_r [2] ? _04216_ : _04213_;
  assign _04218_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [3] : \MSYNC_1r1w.synth.nz.mem[72] [3];
  assign _04219_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [3] : \MSYNC_1r1w.synth.nz.mem[74] [3];
  assign _04220_ = \bapg_rd.w_ptr_r [1] ? _04219_ : _04218_;
  assign _04221_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [3] : \MSYNC_1r1w.synth.nz.mem[76] [3];
  assign _04222_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [3] : \MSYNC_1r1w.synth.nz.mem[78] [3];
  assign _04223_ = \bapg_rd.w_ptr_r [1] ? _04222_ : _04221_;
  assign _04224_ = \bapg_rd.w_ptr_r [2] ? _04223_ : _04220_;
  assign _04225_ = \bapg_rd.w_ptr_r [3] ? _04224_ : _04217_;
  assign _04226_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [3] : \MSYNC_1r1w.synth.nz.mem[80] [3];
  assign _04227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [3] : \MSYNC_1r1w.synth.nz.mem[82] [3];
  assign _04228_ = \bapg_rd.w_ptr_r [1] ? _04227_ : _04226_;
  assign _04229_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [3] : \MSYNC_1r1w.synth.nz.mem[84] [3];
  assign _04230_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [3] : \MSYNC_1r1w.synth.nz.mem[86] [3];
  assign _04231_ = \bapg_rd.w_ptr_r [1] ? _04230_ : _04229_;
  assign _04232_ = \bapg_rd.w_ptr_r [2] ? _04231_ : _04228_;
  assign _04233_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [3] : \MSYNC_1r1w.synth.nz.mem[88] [3];
  assign _04234_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [3] : \MSYNC_1r1w.synth.nz.mem[90] [3];
  assign _04235_ = \bapg_rd.w_ptr_r [1] ? _04234_ : _04233_;
  assign _04236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [3] : \MSYNC_1r1w.synth.nz.mem[92] [3];
  assign _04237_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [3] : \MSYNC_1r1w.synth.nz.mem[94] [3];
  assign _04238_ = \bapg_rd.w_ptr_r [1] ? _04237_ : _04236_;
  assign _04239_ = \bapg_rd.w_ptr_r [2] ? _04238_ : _04235_;
  assign _04240_ = \bapg_rd.w_ptr_r [3] ? _04239_ : _04232_;
  assign _04241_ = \bapg_rd.w_ptr_r [4] ? _04240_ : _04225_;
  assign _04242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [3] : \MSYNC_1r1w.synth.nz.mem[96] [3];
  assign _04243_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [3] : \MSYNC_1r1w.synth.nz.mem[98] [3];
  assign _04244_ = \bapg_rd.w_ptr_r [1] ? _04243_ : _04242_;
  assign _04245_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [3] : \MSYNC_1r1w.synth.nz.mem[100] [3];
  assign _04246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [3] : \MSYNC_1r1w.synth.nz.mem[102] [3];
  assign _04247_ = \bapg_rd.w_ptr_r [1] ? _04246_ : _04245_;
  assign _04248_ = \bapg_rd.w_ptr_r [2] ? _04247_ : _04244_;
  assign _04249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [3] : \MSYNC_1r1w.synth.nz.mem[104] [3];
  assign _04250_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [3] : \MSYNC_1r1w.synth.nz.mem[106] [3];
  assign _04251_ = \bapg_rd.w_ptr_r [1] ? _04250_ : _04249_;
  assign _04252_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [3] : \MSYNC_1r1w.synth.nz.mem[108] [3];
  assign _04253_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [3] : \MSYNC_1r1w.synth.nz.mem[110] [3];
  assign _04254_ = \bapg_rd.w_ptr_r [1] ? _04253_ : _04252_;
  assign _04255_ = \bapg_rd.w_ptr_r [2] ? _04254_ : _04251_;
  assign _04256_ = \bapg_rd.w_ptr_r [3] ? _04255_ : _04248_;
  assign _04257_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [3] : \MSYNC_1r1w.synth.nz.mem[112] [3];
  assign _04258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [3] : \MSYNC_1r1w.synth.nz.mem[114] [3];
  assign _04259_ = \bapg_rd.w_ptr_r [1] ? _04258_ : _04257_;
  assign _04260_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [3] : \MSYNC_1r1w.synth.nz.mem[116] [3];
  assign _04261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [3] : \MSYNC_1r1w.synth.nz.mem[118] [3];
  assign _04262_ = \bapg_rd.w_ptr_r [1] ? _04261_ : _04260_;
  assign _04263_ = \bapg_rd.w_ptr_r [2] ? _04262_ : _04259_;
  assign _04264_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [3] : \MSYNC_1r1w.synth.nz.mem[120] [3];
  assign _04265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [3] : \MSYNC_1r1w.synth.nz.mem[122] [3];
  assign _04266_ = \bapg_rd.w_ptr_r [1] ? _04265_ : _04264_;
  assign _04267_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [3] : \MSYNC_1r1w.synth.nz.mem[124] [3];
  assign _04268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [3] : \MSYNC_1r1w.synth.nz.mem[126] [3];
  assign _04269_ = \bapg_rd.w_ptr_r [1] ? _04268_ : _04267_;
  assign _04270_ = \bapg_rd.w_ptr_r [2] ? _04269_ : _04266_;
  assign _04271_ = \bapg_rd.w_ptr_r [3] ? _04270_ : _04263_;
  assign _04272_ = \bapg_rd.w_ptr_r [4] ? _04271_ : _04256_;
  assign _04273_ = \bapg_rd.w_ptr_r [5] ? _04272_ : _04241_;
  assign _04274_ = \bapg_rd.w_ptr_r [6] ? _04273_ : _04210_;
  assign _04275_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [3] : \MSYNC_1r1w.synth.nz.mem[128] [3];
  assign _04276_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [3] : \MSYNC_1r1w.synth.nz.mem[130] [3];
  assign _04277_ = \bapg_rd.w_ptr_r [1] ? _04276_ : _04275_;
  assign _04278_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [3] : \MSYNC_1r1w.synth.nz.mem[132] [3];
  assign _04279_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [3] : \MSYNC_1r1w.synth.nz.mem[134] [3];
  assign _04280_ = \bapg_rd.w_ptr_r [1] ? _04279_ : _04278_;
  assign _04281_ = \bapg_rd.w_ptr_r [2] ? _04280_ : _04277_;
  assign _04282_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [3] : \MSYNC_1r1w.synth.nz.mem[136] [3];
  assign _04283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [3] : \MSYNC_1r1w.synth.nz.mem[138] [3];
  assign _04284_ = \bapg_rd.w_ptr_r [1] ? _04283_ : _04282_;
  assign _04285_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [3] : \MSYNC_1r1w.synth.nz.mem[140] [3];
  assign _04286_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [3] : \MSYNC_1r1w.synth.nz.mem[142] [3];
  assign _04287_ = \bapg_rd.w_ptr_r [1] ? _04286_ : _04285_;
  assign _04288_ = \bapg_rd.w_ptr_r [2] ? _04287_ : _04284_;
  assign _04289_ = \bapg_rd.w_ptr_r [3] ? _04288_ : _04281_;
  assign _04290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [3] : \MSYNC_1r1w.synth.nz.mem[144] [3];
  assign _04291_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [3] : \MSYNC_1r1w.synth.nz.mem[146] [3];
  assign _04292_ = \bapg_rd.w_ptr_r [1] ? _04291_ : _04290_;
  assign _04293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [3] : \MSYNC_1r1w.synth.nz.mem[148] [3];
  assign _04294_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [3] : \MSYNC_1r1w.synth.nz.mem[150] [3];
  assign _04295_ = \bapg_rd.w_ptr_r [1] ? _04294_ : _04293_;
  assign _04296_ = \bapg_rd.w_ptr_r [2] ? _04295_ : _04292_;
  assign _04297_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [3] : \MSYNC_1r1w.synth.nz.mem[152] [3];
  assign _04298_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [3] : \MSYNC_1r1w.synth.nz.mem[154] [3];
  assign _04299_ = \bapg_rd.w_ptr_r [1] ? _04298_ : _04297_;
  assign _04300_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [3] : \MSYNC_1r1w.synth.nz.mem[156] [3];
  assign _04301_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [3] : \MSYNC_1r1w.synth.nz.mem[158] [3];
  assign _04302_ = \bapg_rd.w_ptr_r [1] ? _04301_ : _04300_;
  assign _04303_ = \bapg_rd.w_ptr_r [2] ? _04302_ : _04299_;
  assign _04304_ = \bapg_rd.w_ptr_r [3] ? _04303_ : _04296_;
  assign _04305_ = \bapg_rd.w_ptr_r [4] ? _04304_ : _04289_;
  assign _04306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [3] : \MSYNC_1r1w.synth.nz.mem[160] [3];
  assign _04307_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [3] : \MSYNC_1r1w.synth.nz.mem[162] [3];
  assign _04308_ = \bapg_rd.w_ptr_r [1] ? _04307_ : _04306_;
  assign _04309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [3] : \MSYNC_1r1w.synth.nz.mem[164] [3];
  assign _04310_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [3] : \MSYNC_1r1w.synth.nz.mem[166] [3];
  assign _04311_ = \bapg_rd.w_ptr_r [1] ? _04310_ : _04309_;
  assign _04312_ = \bapg_rd.w_ptr_r [2] ? _04311_ : _04308_;
  assign _04313_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [3] : \MSYNC_1r1w.synth.nz.mem[168] [3];
  assign _04314_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [3] : \MSYNC_1r1w.synth.nz.mem[170] [3];
  assign _04315_ = \bapg_rd.w_ptr_r [1] ? _04314_ : _04313_;
  assign _04316_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [3] : \MSYNC_1r1w.synth.nz.mem[172] [3];
  assign _04317_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [3] : \MSYNC_1r1w.synth.nz.mem[174] [3];
  assign _04318_ = \bapg_rd.w_ptr_r [1] ? _04317_ : _04316_;
  assign _04319_ = \bapg_rd.w_ptr_r [2] ? _04318_ : _04315_;
  assign _04320_ = \bapg_rd.w_ptr_r [3] ? _04319_ : _04312_;
  assign _04321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [3] : \MSYNC_1r1w.synth.nz.mem[176] [3];
  assign _04322_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [3] : \MSYNC_1r1w.synth.nz.mem[178] [3];
  assign _04323_ = \bapg_rd.w_ptr_r [1] ? _04322_ : _04321_;
  assign _04324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [3] : \MSYNC_1r1w.synth.nz.mem[180] [3];
  assign _04325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [3] : \MSYNC_1r1w.synth.nz.mem[182] [3];
  assign _04326_ = \bapg_rd.w_ptr_r [1] ? _04325_ : _04324_;
  assign _04327_ = \bapg_rd.w_ptr_r [2] ? _04326_ : _04323_;
  assign _04328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [3] : \MSYNC_1r1w.synth.nz.mem[184] [3];
  assign _04329_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [3] : \MSYNC_1r1w.synth.nz.mem[186] [3];
  assign _04330_ = \bapg_rd.w_ptr_r [1] ? _04329_ : _04328_;
  assign _04331_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [3] : \MSYNC_1r1w.synth.nz.mem[188] [3];
  assign _04332_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [3] : \MSYNC_1r1w.synth.nz.mem[190] [3];
  assign _04333_ = \bapg_rd.w_ptr_r [1] ? _04332_ : _04331_;
  assign _04334_ = \bapg_rd.w_ptr_r [2] ? _04333_ : _04330_;
  assign _04335_ = \bapg_rd.w_ptr_r [3] ? _04334_ : _04327_;
  assign _04336_ = \bapg_rd.w_ptr_r [4] ? _04335_ : _04320_;
  assign _04337_ = \bapg_rd.w_ptr_r [5] ? _04336_ : _04305_;
  assign _04338_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [3] : \MSYNC_1r1w.synth.nz.mem[192] [3];
  assign _04339_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [3] : \MSYNC_1r1w.synth.nz.mem[194] [3];
  assign _04340_ = \bapg_rd.w_ptr_r [1] ? _04339_ : _04338_;
  assign _04341_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [3] : \MSYNC_1r1w.synth.nz.mem[196] [3];
  assign _04342_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [3] : \MSYNC_1r1w.synth.nz.mem[198] [3];
  assign _04343_ = \bapg_rd.w_ptr_r [1] ? _04342_ : _04341_;
  assign _04344_ = \bapg_rd.w_ptr_r [2] ? _04343_ : _04340_;
  assign _04345_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [3] : \MSYNC_1r1w.synth.nz.mem[200] [3];
  assign _04346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [3] : \MSYNC_1r1w.synth.nz.mem[202] [3];
  assign _04347_ = \bapg_rd.w_ptr_r [1] ? _04346_ : _04345_;
  assign _04348_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [3] : \MSYNC_1r1w.synth.nz.mem[204] [3];
  assign _04349_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [3] : \MSYNC_1r1w.synth.nz.mem[206] [3];
  assign _04350_ = \bapg_rd.w_ptr_r [1] ? _04349_ : _04348_;
  assign _04351_ = \bapg_rd.w_ptr_r [2] ? _04350_ : _04347_;
  assign _04352_ = \bapg_rd.w_ptr_r [3] ? _04351_ : _04344_;
  assign _04353_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [3] : \MSYNC_1r1w.synth.nz.mem[208] [3];
  assign _04354_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [3] : \MSYNC_1r1w.synth.nz.mem[210] [3];
  assign _04355_ = \bapg_rd.w_ptr_r [1] ? _04354_ : _04353_;
  assign _04356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [3] : \MSYNC_1r1w.synth.nz.mem[212] [3];
  assign _04357_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [3] : \MSYNC_1r1w.synth.nz.mem[214] [3];
  assign _04358_ = \bapg_rd.w_ptr_r [1] ? _04357_ : _04356_;
  assign _04359_ = \bapg_rd.w_ptr_r [2] ? _04358_ : _04355_;
  assign _04360_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [3] : \MSYNC_1r1w.synth.nz.mem[216] [3];
  assign _04361_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [3] : \MSYNC_1r1w.synth.nz.mem[218] [3];
  assign _04362_ = \bapg_rd.w_ptr_r [1] ? _04361_ : _04360_;
  assign _04363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [3] : \MSYNC_1r1w.synth.nz.mem[220] [3];
  assign _04364_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [3] : \MSYNC_1r1w.synth.nz.mem[222] [3];
  assign _04365_ = \bapg_rd.w_ptr_r [1] ? _04364_ : _04363_;
  assign _04366_ = \bapg_rd.w_ptr_r [2] ? _04365_ : _04362_;
  assign _04367_ = \bapg_rd.w_ptr_r [3] ? _04366_ : _04359_;
  assign _04368_ = \bapg_rd.w_ptr_r [4] ? _04367_ : _04352_;
  assign _04369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [3] : \MSYNC_1r1w.synth.nz.mem[224] [3];
  assign _04370_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [3] : \MSYNC_1r1w.synth.nz.mem[226] [3];
  assign _04371_ = \bapg_rd.w_ptr_r [1] ? _04370_ : _04369_;
  assign _04372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [3] : \MSYNC_1r1w.synth.nz.mem[228] [3];
  assign _04373_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [3] : \MSYNC_1r1w.synth.nz.mem[230] [3];
  assign _04374_ = \bapg_rd.w_ptr_r [1] ? _04373_ : _04372_;
  assign _04375_ = \bapg_rd.w_ptr_r [2] ? _04374_ : _04371_;
  assign _04376_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [3] : \MSYNC_1r1w.synth.nz.mem[232] [3];
  assign _04377_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [3] : \MSYNC_1r1w.synth.nz.mem[234] [3];
  assign _04378_ = \bapg_rd.w_ptr_r [1] ? _04377_ : _04376_;
  assign _04379_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [3] : \MSYNC_1r1w.synth.nz.mem[236] [3];
  assign _04380_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [3] : \MSYNC_1r1w.synth.nz.mem[238] [3];
  assign _04381_ = \bapg_rd.w_ptr_r [1] ? _04380_ : _04379_;
  assign _04382_ = \bapg_rd.w_ptr_r [2] ? _04381_ : _04378_;
  assign _04383_ = \bapg_rd.w_ptr_r [3] ? _04382_ : _04375_;
  assign _04384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [3] : \MSYNC_1r1w.synth.nz.mem[240] [3];
  assign _04385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [3] : \MSYNC_1r1w.synth.nz.mem[242] [3];
  assign _04386_ = \bapg_rd.w_ptr_r [1] ? _04385_ : _04384_;
  assign _04387_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [3] : \MSYNC_1r1w.synth.nz.mem[244] [3];
  assign _04388_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [3] : \MSYNC_1r1w.synth.nz.mem[246] [3];
  assign _04389_ = \bapg_rd.w_ptr_r [1] ? _04388_ : _04387_;
  assign _04390_ = \bapg_rd.w_ptr_r [2] ? _04389_ : _04386_;
  assign _04391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [3] : \MSYNC_1r1w.synth.nz.mem[248] [3];
  assign _04392_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [3] : \MSYNC_1r1w.synth.nz.mem[250] [3];
  assign _04393_ = \bapg_rd.w_ptr_r [1] ? _04392_ : _04391_;
  assign _04394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [3] : \MSYNC_1r1w.synth.nz.mem[252] [3];
  assign _04395_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [3] : \MSYNC_1r1w.synth.nz.mem[254] [3];
  assign _04396_ = \bapg_rd.w_ptr_r [1] ? _04395_ : _04394_;
  assign _04397_ = \bapg_rd.w_ptr_r [2] ? _04396_ : _04393_;
  assign _04398_ = \bapg_rd.w_ptr_r [3] ? _04397_ : _04390_;
  assign _04399_ = \bapg_rd.w_ptr_r [4] ? _04398_ : _04383_;
  assign _04400_ = \bapg_rd.w_ptr_r [5] ? _04399_ : _04368_;
  assign _04401_ = \bapg_rd.w_ptr_r [6] ? _04400_ : _04337_;
  assign _04402_ = \bapg_rd.w_ptr_r [7] ? _04401_ : _04274_;
  assign _04403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [3] : \MSYNC_1r1w.synth.nz.mem[256] [3];
  assign _04404_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [3] : \MSYNC_1r1w.synth.nz.mem[258] [3];
  assign _04405_ = \bapg_rd.w_ptr_r [1] ? _04404_ : _04403_;
  assign _04406_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [3] : \MSYNC_1r1w.synth.nz.mem[260] [3];
  assign _04407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [3] : \MSYNC_1r1w.synth.nz.mem[262] [3];
  assign _04408_ = \bapg_rd.w_ptr_r [1] ? _04407_ : _04406_;
  assign _04409_ = \bapg_rd.w_ptr_r [2] ? _04408_ : _04405_;
  assign _04410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [3] : \MSYNC_1r1w.synth.nz.mem[264] [3];
  assign _04411_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [3] : \MSYNC_1r1w.synth.nz.mem[266] [3];
  assign _04412_ = \bapg_rd.w_ptr_r [1] ? _04411_ : _04410_;
  assign _04413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [3] : \MSYNC_1r1w.synth.nz.mem[268] [3];
  assign _04414_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [3] : \MSYNC_1r1w.synth.nz.mem[270] [3];
  assign _04415_ = \bapg_rd.w_ptr_r [1] ? _04414_ : _04413_;
  assign _04416_ = \bapg_rd.w_ptr_r [2] ? _04415_ : _04412_;
  assign _04417_ = \bapg_rd.w_ptr_r [3] ? _04416_ : _04409_;
  assign _04418_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [3] : \MSYNC_1r1w.synth.nz.mem[272] [3];
  assign _04419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [3] : \MSYNC_1r1w.synth.nz.mem[274] [3];
  assign _04420_ = \bapg_rd.w_ptr_r [1] ? _04419_ : _04418_;
  assign _04421_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [3] : \MSYNC_1r1w.synth.nz.mem[276] [3];
  assign _04422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [3] : \MSYNC_1r1w.synth.nz.mem[278] [3];
  assign _04423_ = \bapg_rd.w_ptr_r [1] ? _04422_ : _04421_;
  assign _04424_ = \bapg_rd.w_ptr_r [2] ? _04423_ : _04420_;
  assign _04425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [3] : \MSYNC_1r1w.synth.nz.mem[280] [3];
  assign _04426_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [3] : \MSYNC_1r1w.synth.nz.mem[282] [3];
  assign _04427_ = \bapg_rd.w_ptr_r [1] ? _04426_ : _04425_;
  assign _04428_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [3] : \MSYNC_1r1w.synth.nz.mem[284] [3];
  assign _04429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [3] : \MSYNC_1r1w.synth.nz.mem[286] [3];
  assign _04430_ = \bapg_rd.w_ptr_r [1] ? _04429_ : _04428_;
  assign _04431_ = \bapg_rd.w_ptr_r [2] ? _04430_ : _04427_;
  assign _04432_ = \bapg_rd.w_ptr_r [3] ? _04431_ : _04424_;
  assign _04433_ = \bapg_rd.w_ptr_r [4] ? _04432_ : _04417_;
  assign _04434_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [3] : \MSYNC_1r1w.synth.nz.mem[288] [3];
  assign _04435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [3] : \MSYNC_1r1w.synth.nz.mem[290] [3];
  assign _04436_ = \bapg_rd.w_ptr_r [1] ? _04435_ : _04434_;
  assign _04437_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [3] : \MSYNC_1r1w.synth.nz.mem[292] [3];
  assign _04438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [3] : \MSYNC_1r1w.synth.nz.mem[294] [3];
  assign _04439_ = \bapg_rd.w_ptr_r [1] ? _04438_ : _04437_;
  assign _04440_ = \bapg_rd.w_ptr_r [2] ? _04439_ : _04436_;
  assign _04441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [3] : \MSYNC_1r1w.synth.nz.mem[296] [3];
  assign _04442_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [3] : \MSYNC_1r1w.synth.nz.mem[298] [3];
  assign _04443_ = \bapg_rd.w_ptr_r [1] ? _04442_ : _04441_;
  assign _04444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [3] : \MSYNC_1r1w.synth.nz.mem[300] [3];
  assign _04445_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [3] : \MSYNC_1r1w.synth.nz.mem[302] [3];
  assign _04446_ = \bapg_rd.w_ptr_r [1] ? _04445_ : _04444_;
  assign _04447_ = \bapg_rd.w_ptr_r [2] ? _04446_ : _04443_;
  assign _04448_ = \bapg_rd.w_ptr_r [3] ? _04447_ : _04440_;
  assign _04449_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [3] : \MSYNC_1r1w.synth.nz.mem[304] [3];
  assign _04450_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [3] : \MSYNC_1r1w.synth.nz.mem[306] [3];
  assign _04451_ = \bapg_rd.w_ptr_r [1] ? _04450_ : _04449_;
  assign _04452_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [3] : \MSYNC_1r1w.synth.nz.mem[308] [3];
  assign _04453_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [3] : \MSYNC_1r1w.synth.nz.mem[310] [3];
  assign _04454_ = \bapg_rd.w_ptr_r [1] ? _04453_ : _04452_;
  assign _04455_ = \bapg_rd.w_ptr_r [2] ? _04454_ : _04451_;
  assign _04456_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [3] : \MSYNC_1r1w.synth.nz.mem[312] [3];
  assign _04457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [3] : \MSYNC_1r1w.synth.nz.mem[314] [3];
  assign _04458_ = \bapg_rd.w_ptr_r [1] ? _04457_ : _04456_;
  assign _04459_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [3] : \MSYNC_1r1w.synth.nz.mem[316] [3];
  assign _04460_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [3] : \MSYNC_1r1w.synth.nz.mem[318] [3];
  assign _04461_ = \bapg_rd.w_ptr_r [1] ? _04460_ : _04459_;
  assign _04462_ = \bapg_rd.w_ptr_r [2] ? _04461_ : _04458_;
  assign _04463_ = \bapg_rd.w_ptr_r [3] ? _04462_ : _04455_;
  assign _04464_ = \bapg_rd.w_ptr_r [4] ? _04463_ : _04448_;
  assign _04465_ = \bapg_rd.w_ptr_r [5] ? _04464_ : _04433_;
  assign _04466_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [3] : \MSYNC_1r1w.synth.nz.mem[320] [3];
  assign _04467_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [3] : \MSYNC_1r1w.synth.nz.mem[322] [3];
  assign _04468_ = \bapg_rd.w_ptr_r [1] ? _04467_ : _04466_;
  assign _04469_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [3] : \MSYNC_1r1w.synth.nz.mem[324] [3];
  assign _04470_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [3] : \MSYNC_1r1w.synth.nz.mem[326] [3];
  assign _04471_ = \bapg_rd.w_ptr_r [1] ? _04470_ : _04469_;
  assign _04472_ = \bapg_rd.w_ptr_r [2] ? _04471_ : _04468_;
  assign _04473_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [3] : \MSYNC_1r1w.synth.nz.mem[328] [3];
  assign _04474_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [3] : \MSYNC_1r1w.synth.nz.mem[330] [3];
  assign _04475_ = \bapg_rd.w_ptr_r [1] ? _04474_ : _04473_;
  assign _04476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [3] : \MSYNC_1r1w.synth.nz.mem[332] [3];
  assign _04477_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [3] : \MSYNC_1r1w.synth.nz.mem[334] [3];
  assign _04478_ = \bapg_rd.w_ptr_r [1] ? _04477_ : _04476_;
  assign _04479_ = \bapg_rd.w_ptr_r [2] ? _04478_ : _04475_;
  assign _04480_ = \bapg_rd.w_ptr_r [3] ? _04479_ : _04472_;
  assign _04481_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [3] : \MSYNC_1r1w.synth.nz.mem[336] [3];
  assign _04482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [3] : \MSYNC_1r1w.synth.nz.mem[338] [3];
  assign _04483_ = \bapg_rd.w_ptr_r [1] ? _04482_ : _04481_;
  assign _04484_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [3] : \MSYNC_1r1w.synth.nz.mem[340] [3];
  assign _04485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [3] : \MSYNC_1r1w.synth.nz.mem[342] [3];
  assign _04486_ = \bapg_rd.w_ptr_r [1] ? _04485_ : _04484_;
  assign _04487_ = \bapg_rd.w_ptr_r [2] ? _04486_ : _04483_;
  assign _04488_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [3] : \MSYNC_1r1w.synth.nz.mem[344] [3];
  assign _04489_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [3] : \MSYNC_1r1w.synth.nz.mem[346] [3];
  assign _04490_ = \bapg_rd.w_ptr_r [1] ? _04489_ : _04488_;
  assign _04491_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [3] : \MSYNC_1r1w.synth.nz.mem[348] [3];
  assign _04492_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [3] : \MSYNC_1r1w.synth.nz.mem[350] [3];
  assign _04493_ = \bapg_rd.w_ptr_r [1] ? _04492_ : _04491_;
  assign _04494_ = \bapg_rd.w_ptr_r [2] ? _04493_ : _04490_;
  assign _04495_ = \bapg_rd.w_ptr_r [3] ? _04494_ : _04487_;
  assign _04496_ = \bapg_rd.w_ptr_r [4] ? _04495_ : _04480_;
  assign _04497_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [3] : \MSYNC_1r1w.synth.nz.mem[352] [3];
  assign _04498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [3] : \MSYNC_1r1w.synth.nz.mem[354] [3];
  assign _04499_ = \bapg_rd.w_ptr_r [1] ? _04498_ : _04497_;
  assign _04500_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [3] : \MSYNC_1r1w.synth.nz.mem[356] [3];
  assign _04501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [3] : \MSYNC_1r1w.synth.nz.mem[358] [3];
  assign _04502_ = \bapg_rd.w_ptr_r [1] ? _04501_ : _04500_;
  assign _04503_ = \bapg_rd.w_ptr_r [2] ? _04502_ : _04499_;
  assign _04504_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [3] : \MSYNC_1r1w.synth.nz.mem[360] [3];
  assign _04505_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [3] : \MSYNC_1r1w.synth.nz.mem[362] [3];
  assign _04506_ = \bapg_rd.w_ptr_r [1] ? _04505_ : _04504_;
  assign _04507_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [3] : \MSYNC_1r1w.synth.nz.mem[364] [3];
  assign _04508_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [3] : \MSYNC_1r1w.synth.nz.mem[366] [3];
  assign _04509_ = \bapg_rd.w_ptr_r [1] ? _04508_ : _04507_;
  assign _04510_ = \bapg_rd.w_ptr_r [2] ? _04509_ : _04506_;
  assign _04511_ = \bapg_rd.w_ptr_r [3] ? _04510_ : _04503_;
  assign _04512_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [3] : \MSYNC_1r1w.synth.nz.mem[368] [3];
  assign _04513_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [3] : \MSYNC_1r1w.synth.nz.mem[370] [3];
  assign _04514_ = \bapg_rd.w_ptr_r [1] ? _04513_ : _04512_;
  assign _04515_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [3] : \MSYNC_1r1w.synth.nz.mem[372] [3];
  assign _04516_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [3] : \MSYNC_1r1w.synth.nz.mem[374] [3];
  assign _04517_ = \bapg_rd.w_ptr_r [1] ? _04516_ : _04515_;
  assign _04518_ = \bapg_rd.w_ptr_r [2] ? _04517_ : _04514_;
  assign _04519_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [3] : \MSYNC_1r1w.synth.nz.mem[376] [3];
  assign _04520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [3] : \MSYNC_1r1w.synth.nz.mem[378] [3];
  assign _04521_ = \bapg_rd.w_ptr_r [1] ? _04520_ : _04519_;
  assign _04522_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [3] : \MSYNC_1r1w.synth.nz.mem[380] [3];
  assign _04523_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [3] : \MSYNC_1r1w.synth.nz.mem[382] [3];
  assign _04524_ = \bapg_rd.w_ptr_r [1] ? _04523_ : _04522_;
  assign _04525_ = \bapg_rd.w_ptr_r [2] ? _04524_ : _04521_;
  assign _04526_ = \bapg_rd.w_ptr_r [3] ? _04525_ : _04518_;
  assign _04527_ = \bapg_rd.w_ptr_r [4] ? _04526_ : _04511_;
  assign _04528_ = \bapg_rd.w_ptr_r [5] ? _04527_ : _04496_;
  assign _04529_ = \bapg_rd.w_ptr_r [6] ? _04528_ : _04465_;
  assign _04530_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [3] : \MSYNC_1r1w.synth.nz.mem[384] [3];
  assign _04531_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [3] : \MSYNC_1r1w.synth.nz.mem[386] [3];
  assign _04532_ = \bapg_rd.w_ptr_r [1] ? _04531_ : _04530_;
  assign _04533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [3] : \MSYNC_1r1w.synth.nz.mem[388] [3];
  assign _04534_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [3] : \MSYNC_1r1w.synth.nz.mem[390] [3];
  assign _04535_ = \bapg_rd.w_ptr_r [1] ? _04534_ : _04533_;
  assign _04536_ = \bapg_rd.w_ptr_r [2] ? _04535_ : _04532_;
  assign _04537_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [3] : \MSYNC_1r1w.synth.nz.mem[392] [3];
  assign _04538_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [3] : \MSYNC_1r1w.synth.nz.mem[394] [3];
  assign _04539_ = \bapg_rd.w_ptr_r [1] ? _04538_ : _04537_;
  assign _04540_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [3] : \MSYNC_1r1w.synth.nz.mem[396] [3];
  assign _04541_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [3] : \MSYNC_1r1w.synth.nz.mem[398] [3];
  assign _04542_ = \bapg_rd.w_ptr_r [1] ? _04541_ : _04540_;
  assign _04543_ = \bapg_rd.w_ptr_r [2] ? _04542_ : _04539_;
  assign _04544_ = \bapg_rd.w_ptr_r [3] ? _04543_ : _04536_;
  assign _04545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [3] : \MSYNC_1r1w.synth.nz.mem[400] [3];
  assign _04546_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [3] : \MSYNC_1r1w.synth.nz.mem[402] [3];
  assign _04547_ = \bapg_rd.w_ptr_r [1] ? _04546_ : _04545_;
  assign _04548_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [3] : \MSYNC_1r1w.synth.nz.mem[404] [3];
  assign _04549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [3] : \MSYNC_1r1w.synth.nz.mem[406] [3];
  assign _04550_ = \bapg_rd.w_ptr_r [1] ? _04549_ : _04548_;
  assign _04551_ = \bapg_rd.w_ptr_r [2] ? _04550_ : _04547_;
  assign _04552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [3] : \MSYNC_1r1w.synth.nz.mem[408] [3];
  assign _04553_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [3] : \MSYNC_1r1w.synth.nz.mem[410] [3];
  assign _04554_ = \bapg_rd.w_ptr_r [1] ? _04553_ : _04552_;
  assign _04555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [3] : \MSYNC_1r1w.synth.nz.mem[412] [3];
  assign _04556_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [3] : \MSYNC_1r1w.synth.nz.mem[414] [3];
  assign _04557_ = \bapg_rd.w_ptr_r [1] ? _04556_ : _04555_;
  assign _04558_ = \bapg_rd.w_ptr_r [2] ? _04557_ : _04554_;
  assign _04559_ = \bapg_rd.w_ptr_r [3] ? _04558_ : _04551_;
  assign _04560_ = \bapg_rd.w_ptr_r [4] ? _04559_ : _04544_;
  assign _04561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [3] : \MSYNC_1r1w.synth.nz.mem[416] [3];
  assign _04562_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [3] : \MSYNC_1r1w.synth.nz.mem[418] [3];
  assign _04563_ = \bapg_rd.w_ptr_r [1] ? _04562_ : _04561_;
  assign _04564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [3] : \MSYNC_1r1w.synth.nz.mem[420] [3];
  assign _04565_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [3] : \MSYNC_1r1w.synth.nz.mem[422] [3];
  assign _04566_ = \bapg_rd.w_ptr_r [1] ? _04565_ : _04564_;
  assign _04567_ = \bapg_rd.w_ptr_r [2] ? _04566_ : _04563_;
  assign _04568_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [3] : \MSYNC_1r1w.synth.nz.mem[424] [3];
  assign _04569_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [3] : \MSYNC_1r1w.synth.nz.mem[426] [3];
  assign _04570_ = \bapg_rd.w_ptr_r [1] ? _04569_ : _04568_;
  assign _04571_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [3] : \MSYNC_1r1w.synth.nz.mem[428] [3];
  assign _04572_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [3] : \MSYNC_1r1w.synth.nz.mem[430] [3];
  assign _04573_ = \bapg_rd.w_ptr_r [1] ? _04572_ : _04571_;
  assign _04574_ = \bapg_rd.w_ptr_r [2] ? _04573_ : _04570_;
  assign _04575_ = \bapg_rd.w_ptr_r [3] ? _04574_ : _04567_;
  assign _04576_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [3] : \MSYNC_1r1w.synth.nz.mem[432] [3];
  assign _04577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [3] : \MSYNC_1r1w.synth.nz.mem[434] [3];
  assign _04578_ = \bapg_rd.w_ptr_r [1] ? _04577_ : _04576_;
  assign _04579_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [3] : \MSYNC_1r1w.synth.nz.mem[436] [3];
  assign _04580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [3] : \MSYNC_1r1w.synth.nz.mem[438] [3];
  assign _04581_ = \bapg_rd.w_ptr_r [1] ? _04580_ : _04579_;
  assign _04582_ = \bapg_rd.w_ptr_r [2] ? _04581_ : _04578_;
  assign _04583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [3] : \MSYNC_1r1w.synth.nz.mem[440] [3];
  assign _04584_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [3] : \MSYNC_1r1w.synth.nz.mem[442] [3];
  assign _04585_ = \bapg_rd.w_ptr_r [1] ? _04584_ : _04583_;
  assign _04586_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [3] : \MSYNC_1r1w.synth.nz.mem[444] [3];
  assign _04587_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [3] : \MSYNC_1r1w.synth.nz.mem[446] [3];
  assign _04588_ = \bapg_rd.w_ptr_r [1] ? _04587_ : _04586_;
  assign _04589_ = \bapg_rd.w_ptr_r [2] ? _04588_ : _04585_;
  assign _04590_ = \bapg_rd.w_ptr_r [3] ? _04589_ : _04582_;
  assign _04591_ = \bapg_rd.w_ptr_r [4] ? _04590_ : _04575_;
  assign _04592_ = \bapg_rd.w_ptr_r [5] ? _04591_ : _04560_;
  assign _04593_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [3] : \MSYNC_1r1w.synth.nz.mem[448] [3];
  assign _04594_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [3] : \MSYNC_1r1w.synth.nz.mem[450] [3];
  assign _04595_ = \bapg_rd.w_ptr_r [1] ? _04594_ : _04593_;
  assign _04596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [3] : \MSYNC_1r1w.synth.nz.mem[452] [3];
  assign _04597_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [3] : \MSYNC_1r1w.synth.nz.mem[454] [3];
  assign _04598_ = \bapg_rd.w_ptr_r [1] ? _04597_ : _04596_;
  assign _04599_ = \bapg_rd.w_ptr_r [2] ? _04598_ : _04595_;
  assign _04600_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [3] : \MSYNC_1r1w.synth.nz.mem[456] [3];
  assign _04601_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [3] : \MSYNC_1r1w.synth.nz.mem[458] [3];
  assign _04602_ = \bapg_rd.w_ptr_r [1] ? _04601_ : _04600_;
  assign _04603_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [3] : \MSYNC_1r1w.synth.nz.mem[460] [3];
  assign _04604_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [3] : \MSYNC_1r1w.synth.nz.mem[462] [3];
  assign _04605_ = \bapg_rd.w_ptr_r [1] ? _04604_ : _04603_;
  assign _04606_ = \bapg_rd.w_ptr_r [2] ? _04605_ : _04602_;
  assign _04607_ = \bapg_rd.w_ptr_r [3] ? _04606_ : _04599_;
  assign _04608_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [3] : \MSYNC_1r1w.synth.nz.mem[464] [3];
  assign _04609_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [3] : \MSYNC_1r1w.synth.nz.mem[466] [3];
  assign _04610_ = \bapg_rd.w_ptr_r [1] ? _04609_ : _04608_;
  assign _04611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [3] : \MSYNC_1r1w.synth.nz.mem[468] [3];
  assign _04612_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [3] : \MSYNC_1r1w.synth.nz.mem[470] [3];
  assign _04613_ = \bapg_rd.w_ptr_r [1] ? _04612_ : _04611_;
  assign _04614_ = \bapg_rd.w_ptr_r [2] ? _04613_ : _04610_;
  assign _04615_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [3] : \MSYNC_1r1w.synth.nz.mem[472] [3];
  assign _04616_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [3] : \MSYNC_1r1w.synth.nz.mem[474] [3];
  assign _04617_ = \bapg_rd.w_ptr_r [1] ? _04616_ : _04615_;
  assign _04618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [3] : \MSYNC_1r1w.synth.nz.mem[476] [3];
  assign _04619_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [3] : \MSYNC_1r1w.synth.nz.mem[478] [3];
  assign _04620_ = \bapg_rd.w_ptr_r [1] ? _04619_ : _04618_;
  assign _04621_ = \bapg_rd.w_ptr_r [2] ? _04620_ : _04617_;
  assign _04622_ = \bapg_rd.w_ptr_r [3] ? _04621_ : _04614_;
  assign _04623_ = \bapg_rd.w_ptr_r [4] ? _04622_ : _04607_;
  assign _04624_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [3] : \MSYNC_1r1w.synth.nz.mem[480] [3];
  assign _04625_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [3] : \MSYNC_1r1w.synth.nz.mem[482] [3];
  assign _04626_ = \bapg_rd.w_ptr_r [1] ? _04625_ : _04624_;
  assign _04627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [3] : \MSYNC_1r1w.synth.nz.mem[484] [3];
  assign _04628_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [3] : \MSYNC_1r1w.synth.nz.mem[486] [3];
  assign _04629_ = \bapg_rd.w_ptr_r [1] ? _04628_ : _04627_;
  assign _04630_ = \bapg_rd.w_ptr_r [2] ? _04629_ : _04626_;
  assign _04631_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [3] : \MSYNC_1r1w.synth.nz.mem[488] [3];
  assign _04632_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [3] : \MSYNC_1r1w.synth.nz.mem[490] [3];
  assign _04633_ = \bapg_rd.w_ptr_r [1] ? _04632_ : _04631_;
  assign _04634_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [3] : \MSYNC_1r1w.synth.nz.mem[492] [3];
  assign _04635_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [3] : \MSYNC_1r1w.synth.nz.mem[494] [3];
  assign _04636_ = \bapg_rd.w_ptr_r [1] ? _04635_ : _04634_;
  assign _04637_ = \bapg_rd.w_ptr_r [2] ? _04636_ : _04633_;
  assign _04638_ = \bapg_rd.w_ptr_r [3] ? _04637_ : _04630_;
  assign _04639_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [3] : \MSYNC_1r1w.synth.nz.mem[496] [3];
  assign _04640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [3] : \MSYNC_1r1w.synth.nz.mem[498] [3];
  assign _04641_ = \bapg_rd.w_ptr_r [1] ? _04640_ : _04639_;
  assign _04642_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [3] : \MSYNC_1r1w.synth.nz.mem[500] [3];
  assign _04643_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [3] : \MSYNC_1r1w.synth.nz.mem[502] [3];
  assign _04644_ = \bapg_rd.w_ptr_r [1] ? _04643_ : _04642_;
  assign _04645_ = \bapg_rd.w_ptr_r [2] ? _04644_ : _04641_;
  assign _04646_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [3] : \MSYNC_1r1w.synth.nz.mem[504] [3];
  assign _04647_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [3] : \MSYNC_1r1w.synth.nz.mem[506] [3];
  assign _04648_ = \bapg_rd.w_ptr_r [1] ? _04647_ : _04646_;
  assign _04649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [3] : \MSYNC_1r1w.synth.nz.mem[508] [3];
  assign _04650_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [3] : \MSYNC_1r1w.synth.nz.mem[510] [3];
  assign _04651_ = \bapg_rd.w_ptr_r [1] ? _04650_ : _04649_;
  assign _04652_ = \bapg_rd.w_ptr_r [2] ? _04651_ : _04648_;
  assign _04653_ = \bapg_rd.w_ptr_r [3] ? _04652_ : _04645_;
  assign _04654_ = \bapg_rd.w_ptr_r [4] ? _04653_ : _04638_;
  assign _04655_ = \bapg_rd.w_ptr_r [5] ? _04654_ : _04623_;
  assign _04656_ = \bapg_rd.w_ptr_r [6] ? _04655_ : _04592_;
  assign _04657_ = \bapg_rd.w_ptr_r [7] ? _04656_ : _04529_;
  assign _04658_ = \bapg_rd.w_ptr_r [8] ? _04657_ : _04402_;
  assign _04659_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [3] : \MSYNC_1r1w.synth.nz.mem[512] [3];
  assign _04660_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [3] : \MSYNC_1r1w.synth.nz.mem[514] [3];
  assign _04661_ = \bapg_rd.w_ptr_r [1] ? _04660_ : _04659_;
  assign _04662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [3] : \MSYNC_1r1w.synth.nz.mem[516] [3];
  assign _04663_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [3] : \MSYNC_1r1w.synth.nz.mem[518] [3];
  assign _04664_ = \bapg_rd.w_ptr_r [1] ? _04663_ : _04662_;
  assign _04665_ = \bapg_rd.w_ptr_r [2] ? _04664_ : _04661_;
  assign _04666_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [3] : \MSYNC_1r1w.synth.nz.mem[520] [3];
  assign _04667_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [3] : \MSYNC_1r1w.synth.nz.mem[522] [3];
  assign _04668_ = \bapg_rd.w_ptr_r [1] ? _04667_ : _04666_;
  assign _04669_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [3] : \MSYNC_1r1w.synth.nz.mem[524] [3];
  assign _04670_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [3] : \MSYNC_1r1w.synth.nz.mem[526] [3];
  assign _04671_ = \bapg_rd.w_ptr_r [1] ? _04670_ : _04669_;
  assign _04672_ = \bapg_rd.w_ptr_r [2] ? _04671_ : _04668_;
  assign _04673_ = \bapg_rd.w_ptr_r [3] ? _04672_ : _04665_;
  assign _04674_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [3] : \MSYNC_1r1w.synth.nz.mem[528] [3];
  assign _04675_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [3] : \MSYNC_1r1w.synth.nz.mem[530] [3];
  assign _04676_ = \bapg_rd.w_ptr_r [1] ? _04675_ : _04674_;
  assign _04677_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [3] : \MSYNC_1r1w.synth.nz.mem[532] [3];
  assign _04678_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [3] : \MSYNC_1r1w.synth.nz.mem[534] [3];
  assign _04679_ = \bapg_rd.w_ptr_r [1] ? _04678_ : _04677_;
  assign _04680_ = \bapg_rd.w_ptr_r [2] ? _04679_ : _04676_;
  assign _04681_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [3] : \MSYNC_1r1w.synth.nz.mem[536] [3];
  assign _04682_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [3] : \MSYNC_1r1w.synth.nz.mem[538] [3];
  assign _04683_ = \bapg_rd.w_ptr_r [1] ? _04682_ : _04681_;
  assign _04684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [3] : \MSYNC_1r1w.synth.nz.mem[540] [3];
  assign _04685_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [3] : \MSYNC_1r1w.synth.nz.mem[542] [3];
  assign _04686_ = \bapg_rd.w_ptr_r [1] ? _04685_ : _04684_;
  assign _04687_ = \bapg_rd.w_ptr_r [2] ? _04686_ : _04683_;
  assign _04688_ = \bapg_rd.w_ptr_r [3] ? _04687_ : _04680_;
  assign _04689_ = \bapg_rd.w_ptr_r [4] ? _04688_ : _04673_;
  assign _04690_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [3] : \MSYNC_1r1w.synth.nz.mem[544] [3];
  assign _04691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [3] : \MSYNC_1r1w.synth.nz.mem[546] [3];
  assign _04692_ = \bapg_rd.w_ptr_r [1] ? _04691_ : _04690_;
  assign _04693_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [3] : \MSYNC_1r1w.synth.nz.mem[548] [3];
  assign _04694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [3] : \MSYNC_1r1w.synth.nz.mem[550] [3];
  assign _04695_ = \bapg_rd.w_ptr_r [1] ? _04694_ : _04693_;
  assign _04696_ = \bapg_rd.w_ptr_r [2] ? _04695_ : _04692_;
  assign _04697_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [3] : \MSYNC_1r1w.synth.nz.mem[552] [3];
  assign _04698_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [3] : \MSYNC_1r1w.synth.nz.mem[554] [3];
  assign _04699_ = \bapg_rd.w_ptr_r [1] ? _04698_ : _04697_;
  assign _04700_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [3] : \MSYNC_1r1w.synth.nz.mem[556] [3];
  assign _04701_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [3] : \MSYNC_1r1w.synth.nz.mem[558] [3];
  assign _04702_ = \bapg_rd.w_ptr_r [1] ? _04701_ : _04700_;
  assign _04703_ = \bapg_rd.w_ptr_r [2] ? _04702_ : _04699_;
  assign _04704_ = \bapg_rd.w_ptr_r [3] ? _04703_ : _04696_;
  assign _04705_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [3] : \MSYNC_1r1w.synth.nz.mem[560] [3];
  assign _04706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [3] : \MSYNC_1r1w.synth.nz.mem[562] [3];
  assign _04707_ = \bapg_rd.w_ptr_r [1] ? _04706_ : _04705_;
  assign _04708_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [3] : \MSYNC_1r1w.synth.nz.mem[564] [3];
  assign _04709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [3] : \MSYNC_1r1w.synth.nz.mem[566] [3];
  assign _04710_ = \bapg_rd.w_ptr_r [1] ? _04709_ : _04708_;
  assign _04711_ = \bapg_rd.w_ptr_r [2] ? _04710_ : _04707_;
  assign _04712_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [3] : \MSYNC_1r1w.synth.nz.mem[568] [3];
  assign _04713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [3] : \MSYNC_1r1w.synth.nz.mem[570] [3];
  assign _04714_ = \bapg_rd.w_ptr_r [1] ? _04713_ : _04712_;
  assign _04715_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [3] : \MSYNC_1r1w.synth.nz.mem[572] [3];
  assign _04716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [3] : \MSYNC_1r1w.synth.nz.mem[574] [3];
  assign _04717_ = \bapg_rd.w_ptr_r [1] ? _04716_ : _04715_;
  assign _04718_ = \bapg_rd.w_ptr_r [2] ? _04717_ : _04714_;
  assign _04719_ = \bapg_rd.w_ptr_r [3] ? _04718_ : _04711_;
  assign _04720_ = \bapg_rd.w_ptr_r [4] ? _04719_ : _04704_;
  assign _04721_ = \bapg_rd.w_ptr_r [5] ? _04720_ : _04689_;
  assign _04722_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [3] : \MSYNC_1r1w.synth.nz.mem[576] [3];
  assign _04723_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [3] : \MSYNC_1r1w.synth.nz.mem[578] [3];
  assign _04724_ = \bapg_rd.w_ptr_r [1] ? _04723_ : _04722_;
  assign _04725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [3] : \MSYNC_1r1w.synth.nz.mem[580] [3];
  assign _04726_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [3] : \MSYNC_1r1w.synth.nz.mem[582] [3];
  assign _04727_ = \bapg_rd.w_ptr_r [1] ? _04726_ : _04725_;
  assign _04728_ = \bapg_rd.w_ptr_r [2] ? _04727_ : _04724_;
  assign _04729_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [3] : \MSYNC_1r1w.synth.nz.mem[584] [3];
  assign _04730_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [3] : \MSYNC_1r1w.synth.nz.mem[586] [3];
  assign _04731_ = \bapg_rd.w_ptr_r [1] ? _04730_ : _04729_;
  assign _04732_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [3] : \MSYNC_1r1w.synth.nz.mem[588] [3];
  assign _04733_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [3] : \MSYNC_1r1w.synth.nz.mem[590] [3];
  assign _04734_ = \bapg_rd.w_ptr_r [1] ? _04733_ : _04732_;
  assign _04735_ = \bapg_rd.w_ptr_r [2] ? _04734_ : _04731_;
  assign _04736_ = \bapg_rd.w_ptr_r [3] ? _04735_ : _04728_;
  assign _04737_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [3] : \MSYNC_1r1w.synth.nz.mem[592] [3];
  assign _04738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [3] : \MSYNC_1r1w.synth.nz.mem[594] [3];
  assign _04739_ = \bapg_rd.w_ptr_r [1] ? _04738_ : _04737_;
  assign _04740_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [3] : \MSYNC_1r1w.synth.nz.mem[596] [3];
  assign _04741_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [3] : \MSYNC_1r1w.synth.nz.mem[598] [3];
  assign _04742_ = \bapg_rd.w_ptr_r [1] ? _04741_ : _04740_;
  assign _04743_ = \bapg_rd.w_ptr_r [2] ? _04742_ : _04739_;
  assign _04744_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [3] : \MSYNC_1r1w.synth.nz.mem[600] [3];
  assign _04745_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [3] : \MSYNC_1r1w.synth.nz.mem[602] [3];
  assign _04746_ = \bapg_rd.w_ptr_r [1] ? _04745_ : _04744_;
  assign _04747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [3] : \MSYNC_1r1w.synth.nz.mem[604] [3];
  assign _04748_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [3] : \MSYNC_1r1w.synth.nz.mem[606] [3];
  assign _04749_ = \bapg_rd.w_ptr_r [1] ? _04748_ : _04747_;
  assign _04750_ = \bapg_rd.w_ptr_r [2] ? _04749_ : _04746_;
  assign _04751_ = \bapg_rd.w_ptr_r [3] ? _04750_ : _04743_;
  assign _04752_ = \bapg_rd.w_ptr_r [4] ? _04751_ : _04736_;
  assign _04753_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [3] : \MSYNC_1r1w.synth.nz.mem[608] [3];
  assign _04754_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [3] : \MSYNC_1r1w.synth.nz.mem[610] [3];
  assign _04755_ = \bapg_rd.w_ptr_r [1] ? _04754_ : _04753_;
  assign _04756_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [3] : \MSYNC_1r1w.synth.nz.mem[612] [3];
  assign _04757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [3] : \MSYNC_1r1w.synth.nz.mem[614] [3];
  assign _04758_ = \bapg_rd.w_ptr_r [1] ? _04757_ : _04756_;
  assign _04759_ = \bapg_rd.w_ptr_r [2] ? _04758_ : _04755_;
  assign _04760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [3] : \MSYNC_1r1w.synth.nz.mem[616] [3];
  assign _04761_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [3] : \MSYNC_1r1w.synth.nz.mem[618] [3];
  assign _04762_ = \bapg_rd.w_ptr_r [1] ? _04761_ : _04760_;
  assign _04763_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [3] : \MSYNC_1r1w.synth.nz.mem[620] [3];
  assign _04764_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [3] : \MSYNC_1r1w.synth.nz.mem[622] [3];
  assign _04765_ = \bapg_rd.w_ptr_r [1] ? _04764_ : _04763_;
  assign _04766_ = \bapg_rd.w_ptr_r [2] ? _04765_ : _04762_;
  assign _04767_ = \bapg_rd.w_ptr_r [3] ? _04766_ : _04759_;
  assign _04768_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [3] : \MSYNC_1r1w.synth.nz.mem[624] [3];
  assign _04769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [3] : \MSYNC_1r1w.synth.nz.mem[626] [3];
  assign _04770_ = \bapg_rd.w_ptr_r [1] ? _04769_ : _04768_;
  assign _04771_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [3] : \MSYNC_1r1w.synth.nz.mem[628] [3];
  assign _04772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [3] : \MSYNC_1r1w.synth.nz.mem[630] [3];
  assign _04773_ = \bapg_rd.w_ptr_r [1] ? _04772_ : _04771_;
  assign _04774_ = \bapg_rd.w_ptr_r [2] ? _04773_ : _04770_;
  assign _04775_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [3] : \MSYNC_1r1w.synth.nz.mem[632] [3];
  assign _04776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [3] : \MSYNC_1r1w.synth.nz.mem[634] [3];
  assign _04777_ = \bapg_rd.w_ptr_r [1] ? _04776_ : _04775_;
  assign _04778_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [3] : \MSYNC_1r1w.synth.nz.mem[636] [3];
  assign _04779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [3] : \MSYNC_1r1w.synth.nz.mem[638] [3];
  assign _04780_ = \bapg_rd.w_ptr_r [1] ? _04779_ : _04778_;
  assign _04781_ = \bapg_rd.w_ptr_r [2] ? _04780_ : _04777_;
  assign _04782_ = \bapg_rd.w_ptr_r [3] ? _04781_ : _04774_;
  assign _04783_ = \bapg_rd.w_ptr_r [4] ? _04782_ : _04767_;
  assign _04784_ = \bapg_rd.w_ptr_r [5] ? _04783_ : _04752_;
  assign _04785_ = \bapg_rd.w_ptr_r [6] ? _04784_ : _04721_;
  assign _04786_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [3] : \MSYNC_1r1w.synth.nz.mem[640] [3];
  assign _04787_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [3] : \MSYNC_1r1w.synth.nz.mem[642] [3];
  assign _04788_ = \bapg_rd.w_ptr_r [1] ? _04787_ : _04786_;
  assign _04789_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [3] : \MSYNC_1r1w.synth.nz.mem[644] [3];
  assign _04790_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [3] : \MSYNC_1r1w.synth.nz.mem[646] [3];
  assign _04791_ = \bapg_rd.w_ptr_r [1] ? _04790_ : _04789_;
  assign _04792_ = \bapg_rd.w_ptr_r [2] ? _04791_ : _04788_;
  assign _04793_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [3] : \MSYNC_1r1w.synth.nz.mem[648] [3];
  assign _04794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [3] : \MSYNC_1r1w.synth.nz.mem[650] [3];
  assign _04795_ = \bapg_rd.w_ptr_r [1] ? _04794_ : _04793_;
  assign _04796_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [3] : \MSYNC_1r1w.synth.nz.mem[652] [3];
  assign _04797_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [3] : \MSYNC_1r1w.synth.nz.mem[654] [3];
  assign _04798_ = \bapg_rd.w_ptr_r [1] ? _04797_ : _04796_;
  assign _04799_ = \bapg_rd.w_ptr_r [2] ? _04798_ : _04795_;
  assign _04800_ = \bapg_rd.w_ptr_r [3] ? _04799_ : _04792_;
  assign _04801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [3] : \MSYNC_1r1w.synth.nz.mem[656] [3];
  assign _04802_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [3] : \MSYNC_1r1w.synth.nz.mem[658] [3];
  assign _04803_ = \bapg_rd.w_ptr_r [1] ? _04802_ : _04801_;
  assign _04804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [3] : \MSYNC_1r1w.synth.nz.mem[660] [3];
  assign _04805_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [3] : \MSYNC_1r1w.synth.nz.mem[662] [3];
  assign _04806_ = \bapg_rd.w_ptr_r [1] ? _04805_ : _04804_;
  assign _04807_ = \bapg_rd.w_ptr_r [2] ? _04806_ : _04803_;
  assign _04808_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [3] : \MSYNC_1r1w.synth.nz.mem[664] [3];
  assign _04809_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [3] : \MSYNC_1r1w.synth.nz.mem[666] [3];
  assign _04810_ = \bapg_rd.w_ptr_r [1] ? _04809_ : _04808_;
  assign _04811_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [3] : \MSYNC_1r1w.synth.nz.mem[668] [3];
  assign _04812_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [3] : \MSYNC_1r1w.synth.nz.mem[670] [3];
  assign _04813_ = \bapg_rd.w_ptr_r [1] ? _04812_ : _04811_;
  assign _04814_ = \bapg_rd.w_ptr_r [2] ? _04813_ : _04810_;
  assign _04815_ = \bapg_rd.w_ptr_r [3] ? _04814_ : _04807_;
  assign _04816_ = \bapg_rd.w_ptr_r [4] ? _04815_ : _04800_;
  assign _04817_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [3] : \MSYNC_1r1w.synth.nz.mem[672] [3];
  assign _04818_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [3] : \MSYNC_1r1w.synth.nz.mem[674] [3];
  assign _04819_ = \bapg_rd.w_ptr_r [1] ? _04818_ : _04817_;
  assign _04820_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [3] : \MSYNC_1r1w.synth.nz.mem[676] [3];
  assign _04821_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [3] : \MSYNC_1r1w.synth.nz.mem[678] [3];
  assign _04822_ = \bapg_rd.w_ptr_r [1] ? _04821_ : _04820_;
  assign _04823_ = \bapg_rd.w_ptr_r [2] ? _04822_ : _04819_;
  assign _04824_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [3] : \MSYNC_1r1w.synth.nz.mem[680] [3];
  assign _04825_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [3] : \MSYNC_1r1w.synth.nz.mem[682] [3];
  assign _04826_ = \bapg_rd.w_ptr_r [1] ? _04825_ : _04824_;
  assign _04827_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [3] : \MSYNC_1r1w.synth.nz.mem[684] [3];
  assign _04828_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [3] : \MSYNC_1r1w.synth.nz.mem[686] [3];
  assign _04829_ = \bapg_rd.w_ptr_r [1] ? _04828_ : _04827_;
  assign _04830_ = \bapg_rd.w_ptr_r [2] ? _04829_ : _04826_;
  assign _04831_ = \bapg_rd.w_ptr_r [3] ? _04830_ : _04823_;
  assign _04832_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [3] : \MSYNC_1r1w.synth.nz.mem[688] [3];
  assign _04833_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [3] : \MSYNC_1r1w.synth.nz.mem[690] [3];
  assign _04834_ = \bapg_rd.w_ptr_r [1] ? _04833_ : _04832_;
  assign _04835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [3] : \MSYNC_1r1w.synth.nz.mem[692] [3];
  assign _04836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [3] : \MSYNC_1r1w.synth.nz.mem[694] [3];
  assign _04837_ = \bapg_rd.w_ptr_r [1] ? _04836_ : _04835_;
  assign _04838_ = \bapg_rd.w_ptr_r [2] ? _04837_ : _04834_;
  assign _04839_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [3] : \MSYNC_1r1w.synth.nz.mem[696] [3];
  assign _04840_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [3] : \MSYNC_1r1w.synth.nz.mem[698] [3];
  assign _04841_ = \bapg_rd.w_ptr_r [1] ? _04840_ : _04839_;
  assign _04842_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [3] : \MSYNC_1r1w.synth.nz.mem[700] [3];
  assign _04843_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [3] : \MSYNC_1r1w.synth.nz.mem[702] [3];
  assign _04844_ = \bapg_rd.w_ptr_r [1] ? _04843_ : _04842_;
  assign _04845_ = \bapg_rd.w_ptr_r [2] ? _04844_ : _04841_;
  assign _04846_ = \bapg_rd.w_ptr_r [3] ? _04845_ : _04838_;
  assign _04847_ = \bapg_rd.w_ptr_r [4] ? _04846_ : _04831_;
  assign _04848_ = \bapg_rd.w_ptr_r [5] ? _04847_ : _04816_;
  assign _04849_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [3] : \MSYNC_1r1w.synth.nz.mem[704] [3];
  assign _04850_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [3] : \MSYNC_1r1w.synth.nz.mem[706] [3];
  assign _04851_ = \bapg_rd.w_ptr_r [1] ? _04850_ : _04849_;
  assign _04852_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [3] : \MSYNC_1r1w.synth.nz.mem[708] [3];
  assign _04853_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [3] : \MSYNC_1r1w.synth.nz.mem[710] [3];
  assign _04854_ = \bapg_rd.w_ptr_r [1] ? _04853_ : _04852_;
  assign _04855_ = \bapg_rd.w_ptr_r [2] ? _04854_ : _04851_;
  assign _04856_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [3] : \MSYNC_1r1w.synth.nz.mem[712] [3];
  assign _04857_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [3] : \MSYNC_1r1w.synth.nz.mem[714] [3];
  assign _04858_ = \bapg_rd.w_ptr_r [1] ? _04857_ : _04856_;
  assign _04859_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [3] : \MSYNC_1r1w.synth.nz.mem[716] [3];
  assign _04860_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [3] : \MSYNC_1r1w.synth.nz.mem[718] [3];
  assign _04861_ = \bapg_rd.w_ptr_r [1] ? _04860_ : _04859_;
  assign _04862_ = \bapg_rd.w_ptr_r [2] ? _04861_ : _04858_;
  assign _04863_ = \bapg_rd.w_ptr_r [3] ? _04862_ : _04855_;
  assign _04864_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [3] : \MSYNC_1r1w.synth.nz.mem[720] [3];
  assign _04865_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [3] : \MSYNC_1r1w.synth.nz.mem[722] [3];
  assign _04866_ = \bapg_rd.w_ptr_r [1] ? _04865_ : _04864_;
  assign _04867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [3] : \MSYNC_1r1w.synth.nz.mem[724] [3];
  assign _04868_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [3] : \MSYNC_1r1w.synth.nz.mem[726] [3];
  assign _04869_ = \bapg_rd.w_ptr_r [1] ? _04868_ : _04867_;
  assign _04870_ = \bapg_rd.w_ptr_r [2] ? _04869_ : _04866_;
  assign _04871_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [3] : \MSYNC_1r1w.synth.nz.mem[728] [3];
  assign _04872_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [3] : \MSYNC_1r1w.synth.nz.mem[730] [3];
  assign _04873_ = \bapg_rd.w_ptr_r [1] ? _04872_ : _04871_;
  assign _04874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [3] : \MSYNC_1r1w.synth.nz.mem[732] [3];
  assign _04875_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [3] : \MSYNC_1r1w.synth.nz.mem[734] [3];
  assign _04876_ = \bapg_rd.w_ptr_r [1] ? _04875_ : _04874_;
  assign _04877_ = \bapg_rd.w_ptr_r [2] ? _04876_ : _04873_;
  assign _04878_ = \bapg_rd.w_ptr_r [3] ? _04877_ : _04870_;
  assign _04879_ = \bapg_rd.w_ptr_r [4] ? _04878_ : _04863_;
  assign _04880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [3] : \MSYNC_1r1w.synth.nz.mem[736] [3];
  assign _04881_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [3] : \MSYNC_1r1w.synth.nz.mem[738] [3];
  assign _04882_ = \bapg_rd.w_ptr_r [1] ? _04881_ : _04880_;
  assign _04883_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [3] : \MSYNC_1r1w.synth.nz.mem[740] [3];
  assign _04884_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [3] : \MSYNC_1r1w.synth.nz.mem[742] [3];
  assign _04885_ = \bapg_rd.w_ptr_r [1] ? _04884_ : _04883_;
  assign _04886_ = \bapg_rd.w_ptr_r [2] ? _04885_ : _04882_;
  assign _04887_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [3] : \MSYNC_1r1w.synth.nz.mem[744] [3];
  assign _04888_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [3] : \MSYNC_1r1w.synth.nz.mem[746] [3];
  assign _04889_ = \bapg_rd.w_ptr_r [1] ? _04888_ : _04887_;
  assign _04890_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [3] : \MSYNC_1r1w.synth.nz.mem[748] [3];
  assign _04891_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [3] : \MSYNC_1r1w.synth.nz.mem[750] [3];
  assign _04892_ = \bapg_rd.w_ptr_r [1] ? _04891_ : _04890_;
  assign _04893_ = \bapg_rd.w_ptr_r [2] ? _04892_ : _04889_;
  assign _04894_ = \bapg_rd.w_ptr_r [3] ? _04893_ : _04886_;
  assign _04895_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [3] : \MSYNC_1r1w.synth.nz.mem[752] [3];
  assign _04896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [3] : \MSYNC_1r1w.synth.nz.mem[754] [3];
  assign _04897_ = \bapg_rd.w_ptr_r [1] ? _04896_ : _04895_;
  assign _04898_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [3] : \MSYNC_1r1w.synth.nz.mem[756] [3];
  assign _04899_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [3] : \MSYNC_1r1w.synth.nz.mem[758] [3];
  assign _04900_ = \bapg_rd.w_ptr_r [1] ? _04899_ : _04898_;
  assign _04901_ = \bapg_rd.w_ptr_r [2] ? _04900_ : _04897_;
  assign _04902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [3] : \MSYNC_1r1w.synth.nz.mem[760] [3];
  assign _04903_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [3] : \MSYNC_1r1w.synth.nz.mem[762] [3];
  assign _04904_ = \bapg_rd.w_ptr_r [1] ? _04903_ : _04902_;
  assign _04905_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [3] : \MSYNC_1r1w.synth.nz.mem[764] [3];
  assign _04906_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [3] : \MSYNC_1r1w.synth.nz.mem[766] [3];
  assign _04907_ = \bapg_rd.w_ptr_r [1] ? _04906_ : _04905_;
  assign _04908_ = \bapg_rd.w_ptr_r [2] ? _04907_ : _04904_;
  assign _04909_ = \bapg_rd.w_ptr_r [3] ? _04908_ : _04901_;
  assign _04910_ = \bapg_rd.w_ptr_r [4] ? _04909_ : _04894_;
  assign _04911_ = \bapg_rd.w_ptr_r [5] ? _04910_ : _04879_;
  assign _04912_ = \bapg_rd.w_ptr_r [6] ? _04911_ : _04848_;
  assign _04913_ = \bapg_rd.w_ptr_r [7] ? _04912_ : _04785_;
  assign _04914_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [3] : \MSYNC_1r1w.synth.nz.mem[768] [3];
  assign _04915_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [3] : \MSYNC_1r1w.synth.nz.mem[770] [3];
  assign _04916_ = \bapg_rd.w_ptr_r [1] ? _04915_ : _04914_;
  assign _04917_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [3] : \MSYNC_1r1w.synth.nz.mem[772] [3];
  assign _04918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [3] : \MSYNC_1r1w.synth.nz.mem[774] [3];
  assign _04919_ = \bapg_rd.w_ptr_r [1] ? _04918_ : _04917_;
  assign _04920_ = \bapg_rd.w_ptr_r [2] ? _04919_ : _04916_;
  assign _04921_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [3] : \MSYNC_1r1w.synth.nz.mem[776] [3];
  assign _04922_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [3] : \MSYNC_1r1w.synth.nz.mem[778] [3];
  assign _04923_ = \bapg_rd.w_ptr_r [1] ? _04922_ : _04921_;
  assign _04924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [3] : \MSYNC_1r1w.synth.nz.mem[780] [3];
  assign _04925_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [3] : \MSYNC_1r1w.synth.nz.mem[782] [3];
  assign _04926_ = \bapg_rd.w_ptr_r [1] ? _04925_ : _04924_;
  assign _04927_ = \bapg_rd.w_ptr_r [2] ? _04926_ : _04923_;
  assign _04928_ = \bapg_rd.w_ptr_r [3] ? _04927_ : _04920_;
  assign _04929_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [3] : \MSYNC_1r1w.synth.nz.mem[784] [3];
  assign _04930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [3] : \MSYNC_1r1w.synth.nz.mem[786] [3];
  assign _04931_ = \bapg_rd.w_ptr_r [1] ? _04930_ : _04929_;
  assign _04932_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [3] : \MSYNC_1r1w.synth.nz.mem[788] [3];
  assign _04933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [3] : \MSYNC_1r1w.synth.nz.mem[790] [3];
  assign _04934_ = \bapg_rd.w_ptr_r [1] ? _04933_ : _04932_;
  assign _04935_ = \bapg_rd.w_ptr_r [2] ? _04934_ : _04931_;
  assign _04936_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [3] : \MSYNC_1r1w.synth.nz.mem[792] [3];
  assign _04937_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [3] : \MSYNC_1r1w.synth.nz.mem[794] [3];
  assign _04938_ = \bapg_rd.w_ptr_r [1] ? _04937_ : _04936_;
  assign _04939_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [3] : \MSYNC_1r1w.synth.nz.mem[796] [3];
  assign _04940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [3] : \MSYNC_1r1w.synth.nz.mem[798] [3];
  assign _04941_ = \bapg_rd.w_ptr_r [1] ? _04940_ : _04939_;
  assign _04942_ = \bapg_rd.w_ptr_r [2] ? _04941_ : _04938_;
  assign _04943_ = \bapg_rd.w_ptr_r [3] ? _04942_ : _04935_;
  assign _04944_ = \bapg_rd.w_ptr_r [4] ? _04943_ : _04928_;
  assign _04945_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [3] : \MSYNC_1r1w.synth.nz.mem[800] [3];
  assign _04946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [3] : \MSYNC_1r1w.synth.nz.mem[802] [3];
  assign _04947_ = \bapg_rd.w_ptr_r [1] ? _04946_ : _04945_;
  assign _04948_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [3] : \MSYNC_1r1w.synth.nz.mem[804] [3];
  assign _04949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [3] : \MSYNC_1r1w.synth.nz.mem[806] [3];
  assign _04950_ = \bapg_rd.w_ptr_r [1] ? _04949_ : _04948_;
  assign _04951_ = \bapg_rd.w_ptr_r [2] ? _04950_ : _04947_;
  assign _04952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [3] : \MSYNC_1r1w.synth.nz.mem[808] [3];
  assign _04953_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [3] : \MSYNC_1r1w.synth.nz.mem[810] [3];
  assign _04954_ = \bapg_rd.w_ptr_r [1] ? _04953_ : _04952_;
  assign _04955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [3] : \MSYNC_1r1w.synth.nz.mem[812] [3];
  assign _04956_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [3] : \MSYNC_1r1w.synth.nz.mem[814] [3];
  assign _04957_ = \bapg_rd.w_ptr_r [1] ? _04956_ : _04955_;
  assign _04958_ = \bapg_rd.w_ptr_r [2] ? _04957_ : _04954_;
  assign _04959_ = \bapg_rd.w_ptr_r [3] ? _04958_ : _04951_;
  assign _04960_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [3] : \MSYNC_1r1w.synth.nz.mem[816] [3];
  assign _04961_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [3] : \MSYNC_1r1w.synth.nz.mem[818] [3];
  assign _04962_ = \bapg_rd.w_ptr_r [1] ? _04961_ : _04960_;
  assign _04963_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [3] : \MSYNC_1r1w.synth.nz.mem[820] [3];
  assign _04964_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [3] : \MSYNC_1r1w.synth.nz.mem[822] [3];
  assign _04965_ = \bapg_rd.w_ptr_r [1] ? _04964_ : _04963_;
  assign _04966_ = \bapg_rd.w_ptr_r [2] ? _04965_ : _04962_;
  assign _04967_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [3] : \MSYNC_1r1w.synth.nz.mem[824] [3];
  assign _04968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [3] : \MSYNC_1r1w.synth.nz.mem[826] [3];
  assign _04969_ = \bapg_rd.w_ptr_r [1] ? _04968_ : _04967_;
  assign _04970_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [3] : \MSYNC_1r1w.synth.nz.mem[828] [3];
  assign _04971_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [3] : \MSYNC_1r1w.synth.nz.mem[830] [3];
  assign _04972_ = \bapg_rd.w_ptr_r [1] ? _04971_ : _04970_;
  assign _04973_ = \bapg_rd.w_ptr_r [2] ? _04972_ : _04969_;
  assign _04974_ = \bapg_rd.w_ptr_r [3] ? _04973_ : _04966_;
  assign _04975_ = \bapg_rd.w_ptr_r [4] ? _04974_ : _04959_;
  assign _04976_ = \bapg_rd.w_ptr_r [5] ? _04975_ : _04944_;
  assign _04977_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [3] : \MSYNC_1r1w.synth.nz.mem[832] [3];
  assign _04978_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [3] : \MSYNC_1r1w.synth.nz.mem[834] [3];
  assign _04979_ = \bapg_rd.w_ptr_r [1] ? _04978_ : _04977_;
  assign _04980_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [3] : \MSYNC_1r1w.synth.nz.mem[836] [3];
  assign _04981_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [3] : \MSYNC_1r1w.synth.nz.mem[838] [3];
  assign _04982_ = \bapg_rd.w_ptr_r [1] ? _04981_ : _04980_;
  assign _04983_ = \bapg_rd.w_ptr_r [2] ? _04982_ : _04979_;
  assign _04984_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [3] : \MSYNC_1r1w.synth.nz.mem[840] [3];
  assign _04985_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [3] : \MSYNC_1r1w.synth.nz.mem[842] [3];
  assign _04986_ = \bapg_rd.w_ptr_r [1] ? _04985_ : _04984_;
  assign _04987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [3] : \MSYNC_1r1w.synth.nz.mem[844] [3];
  assign _04988_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [3] : \MSYNC_1r1w.synth.nz.mem[846] [3];
  assign _04989_ = \bapg_rd.w_ptr_r [1] ? _04988_ : _04987_;
  assign _04990_ = \bapg_rd.w_ptr_r [2] ? _04989_ : _04986_;
  assign _04991_ = \bapg_rd.w_ptr_r [3] ? _04990_ : _04983_;
  assign _04992_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [3] : \MSYNC_1r1w.synth.nz.mem[848] [3];
  assign _04993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [3] : \MSYNC_1r1w.synth.nz.mem[850] [3];
  assign _04994_ = \bapg_rd.w_ptr_r [1] ? _04993_ : _04992_;
  assign _04995_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [3] : \MSYNC_1r1w.synth.nz.mem[852] [3];
  assign _04996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [3] : \MSYNC_1r1w.synth.nz.mem[854] [3];
  assign _04997_ = \bapg_rd.w_ptr_r [1] ? _04996_ : _04995_;
  assign _04998_ = \bapg_rd.w_ptr_r [2] ? _04997_ : _04994_;
  assign _04999_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [3] : \MSYNC_1r1w.synth.nz.mem[856] [3];
  assign _05000_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [3] : \MSYNC_1r1w.synth.nz.mem[858] [3];
  assign _05001_ = \bapg_rd.w_ptr_r [1] ? _05000_ : _04999_;
  assign _05002_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [3] : \MSYNC_1r1w.synth.nz.mem[860] [3];
  assign _05003_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [3] : \MSYNC_1r1w.synth.nz.mem[862] [3];
  assign _05004_ = \bapg_rd.w_ptr_r [1] ? _05003_ : _05002_;
  assign _05005_ = \bapg_rd.w_ptr_r [2] ? _05004_ : _05001_;
  assign _05006_ = \bapg_rd.w_ptr_r [3] ? _05005_ : _04998_;
  assign _05007_ = \bapg_rd.w_ptr_r [4] ? _05006_ : _04991_;
  assign _05008_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [3] : \MSYNC_1r1w.synth.nz.mem[864] [3];
  assign _05009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [3] : \MSYNC_1r1w.synth.nz.mem[866] [3];
  assign _05010_ = \bapg_rd.w_ptr_r [1] ? _05009_ : _05008_;
  assign _05011_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [3] : \MSYNC_1r1w.synth.nz.mem[868] [3];
  assign _05012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [3] : \MSYNC_1r1w.synth.nz.mem[870] [3];
  assign _05013_ = \bapg_rd.w_ptr_r [1] ? _05012_ : _05011_;
  assign _05014_ = \bapg_rd.w_ptr_r [2] ? _05013_ : _05010_;
  assign _05015_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [3] : \MSYNC_1r1w.synth.nz.mem[872] [3];
  assign _05016_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [3] : \MSYNC_1r1w.synth.nz.mem[874] [3];
  assign _05017_ = \bapg_rd.w_ptr_r [1] ? _05016_ : _05015_;
  assign _05018_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [3] : \MSYNC_1r1w.synth.nz.mem[876] [3];
  assign _05019_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [3] : \MSYNC_1r1w.synth.nz.mem[878] [3];
  assign _05020_ = \bapg_rd.w_ptr_r [1] ? _05019_ : _05018_;
  assign _05021_ = \bapg_rd.w_ptr_r [2] ? _05020_ : _05017_;
  assign _05022_ = \bapg_rd.w_ptr_r [3] ? _05021_ : _05014_;
  assign _05023_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [3] : \MSYNC_1r1w.synth.nz.mem[880] [3];
  assign _05024_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [3] : \MSYNC_1r1w.synth.nz.mem[882] [3];
  assign _05025_ = \bapg_rd.w_ptr_r [1] ? _05024_ : _05023_;
  assign _05026_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [3] : \MSYNC_1r1w.synth.nz.mem[884] [3];
  assign _05027_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [3] : \MSYNC_1r1w.synth.nz.mem[886] [3];
  assign _05028_ = \bapg_rd.w_ptr_r [1] ? _05027_ : _05026_;
  assign _05029_ = \bapg_rd.w_ptr_r [2] ? _05028_ : _05025_;
  assign _05030_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [3] : \MSYNC_1r1w.synth.nz.mem[888] [3];
  assign _05031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [3] : \MSYNC_1r1w.synth.nz.mem[890] [3];
  assign _05032_ = \bapg_rd.w_ptr_r [1] ? _05031_ : _05030_;
  assign _05033_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [3] : \MSYNC_1r1w.synth.nz.mem[892] [3];
  assign _05034_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [3] : \MSYNC_1r1w.synth.nz.mem[894] [3];
  assign _05035_ = \bapg_rd.w_ptr_r [1] ? _05034_ : _05033_;
  assign _05036_ = \bapg_rd.w_ptr_r [2] ? _05035_ : _05032_;
  assign _05037_ = \bapg_rd.w_ptr_r [3] ? _05036_ : _05029_;
  assign _05038_ = \bapg_rd.w_ptr_r [4] ? _05037_ : _05022_;
  assign _05039_ = \bapg_rd.w_ptr_r [5] ? _05038_ : _05007_;
  assign _05040_ = \bapg_rd.w_ptr_r [6] ? _05039_ : _04976_;
  assign _05041_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [3] : \MSYNC_1r1w.synth.nz.mem[896] [3];
  assign _05042_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [3] : \MSYNC_1r1w.synth.nz.mem[898] [3];
  assign _05043_ = \bapg_rd.w_ptr_r [1] ? _05042_ : _05041_;
  assign _05044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [3] : \MSYNC_1r1w.synth.nz.mem[900] [3];
  assign _05045_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [3] : \MSYNC_1r1w.synth.nz.mem[902] [3];
  assign _05046_ = \bapg_rd.w_ptr_r [1] ? _05045_ : _05044_;
  assign _05047_ = \bapg_rd.w_ptr_r [2] ? _05046_ : _05043_;
  assign _05048_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [3] : \MSYNC_1r1w.synth.nz.mem[904] [3];
  assign _05049_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [3] : \MSYNC_1r1w.synth.nz.mem[906] [3];
  assign _05050_ = \bapg_rd.w_ptr_r [1] ? _05049_ : _05048_;
  assign _05051_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [3] : \MSYNC_1r1w.synth.nz.mem[908] [3];
  assign _05052_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [3] : \MSYNC_1r1w.synth.nz.mem[910] [3];
  assign _05053_ = \bapg_rd.w_ptr_r [1] ? _05052_ : _05051_;
  assign _05054_ = \bapg_rd.w_ptr_r [2] ? _05053_ : _05050_;
  assign _05055_ = \bapg_rd.w_ptr_r [3] ? _05054_ : _05047_;
  assign _05056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [3] : \MSYNC_1r1w.synth.nz.mem[912] [3];
  assign _05057_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [3] : \MSYNC_1r1w.synth.nz.mem[914] [3];
  assign _05058_ = \bapg_rd.w_ptr_r [1] ? _05057_ : _05056_;
  assign _05059_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [3] : \MSYNC_1r1w.synth.nz.mem[916] [3];
  assign _05060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [3] : \MSYNC_1r1w.synth.nz.mem[918] [3];
  assign _05061_ = \bapg_rd.w_ptr_r [1] ? _05060_ : _05059_;
  assign _05062_ = \bapg_rd.w_ptr_r [2] ? _05061_ : _05058_;
  assign _05063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [3] : \MSYNC_1r1w.synth.nz.mem[920] [3];
  assign _05064_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [3] : \MSYNC_1r1w.synth.nz.mem[922] [3];
  assign _05065_ = \bapg_rd.w_ptr_r [1] ? _05064_ : _05063_;
  assign _05066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [3] : \MSYNC_1r1w.synth.nz.mem[924] [3];
  assign _05067_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [3] : \MSYNC_1r1w.synth.nz.mem[926] [3];
  assign _05068_ = \bapg_rd.w_ptr_r [1] ? _05067_ : _05066_;
  assign _05069_ = \bapg_rd.w_ptr_r [2] ? _05068_ : _05065_;
  assign _05070_ = \bapg_rd.w_ptr_r [3] ? _05069_ : _05062_;
  assign _05071_ = \bapg_rd.w_ptr_r [4] ? _05070_ : _05055_;
  assign _05072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [3] : \MSYNC_1r1w.synth.nz.mem[928] [3];
  assign _05073_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [3] : \MSYNC_1r1w.synth.nz.mem[930] [3];
  assign _05074_ = \bapg_rd.w_ptr_r [1] ? _05073_ : _05072_;
  assign _05075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [3] : \MSYNC_1r1w.synth.nz.mem[932] [3];
  assign _05076_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [3] : \MSYNC_1r1w.synth.nz.mem[934] [3];
  assign _05077_ = \bapg_rd.w_ptr_r [1] ? _05076_ : _05075_;
  assign _05078_ = \bapg_rd.w_ptr_r [2] ? _05077_ : _05074_;
  assign _05079_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [3] : \MSYNC_1r1w.synth.nz.mem[936] [3];
  assign _05080_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [3] : \MSYNC_1r1w.synth.nz.mem[938] [3];
  assign _05081_ = \bapg_rd.w_ptr_r [1] ? _05080_ : _05079_;
  assign _05082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [3] : \MSYNC_1r1w.synth.nz.mem[940] [3];
  assign _05083_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [3] : \MSYNC_1r1w.synth.nz.mem[942] [3];
  assign _05084_ = \bapg_rd.w_ptr_r [1] ? _05083_ : _05082_;
  assign _05085_ = \bapg_rd.w_ptr_r [2] ? _05084_ : _05081_;
  assign _05086_ = \bapg_rd.w_ptr_r [3] ? _05085_ : _05078_;
  assign _05087_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [3] : \MSYNC_1r1w.synth.nz.mem[944] [3];
  assign _05088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [3] : \MSYNC_1r1w.synth.nz.mem[946] [3];
  assign _05089_ = \bapg_rd.w_ptr_r [1] ? _05088_ : _05087_;
  assign _05090_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [3] : \MSYNC_1r1w.synth.nz.mem[948] [3];
  assign _05091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [3] : \MSYNC_1r1w.synth.nz.mem[950] [3];
  assign _05092_ = \bapg_rd.w_ptr_r [1] ? _05091_ : _05090_;
  assign _05093_ = \bapg_rd.w_ptr_r [2] ? _05092_ : _05089_;
  assign _05094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [3] : \MSYNC_1r1w.synth.nz.mem[952] [3];
  assign _05095_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [3] : \MSYNC_1r1w.synth.nz.mem[954] [3];
  assign _05096_ = \bapg_rd.w_ptr_r [1] ? _05095_ : _05094_;
  assign _05097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [3] : \MSYNC_1r1w.synth.nz.mem[956] [3];
  assign _05098_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [3] : \MSYNC_1r1w.synth.nz.mem[958] [3];
  assign _05099_ = \bapg_rd.w_ptr_r [1] ? _05098_ : _05097_;
  assign _05100_ = \bapg_rd.w_ptr_r [2] ? _05099_ : _05096_;
  assign _05101_ = \bapg_rd.w_ptr_r [3] ? _05100_ : _05093_;
  assign _05102_ = \bapg_rd.w_ptr_r [4] ? _05101_ : _05086_;
  assign _05103_ = \bapg_rd.w_ptr_r [5] ? _05102_ : _05071_;
  assign _05104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [3] : \MSYNC_1r1w.synth.nz.mem[960] [3];
  assign _05105_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [3] : \MSYNC_1r1w.synth.nz.mem[962] [3];
  assign _05106_ = \bapg_rd.w_ptr_r [1] ? _05105_ : _05104_;
  assign _05107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [3] : \MSYNC_1r1w.synth.nz.mem[964] [3];
  assign _05108_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [3] : \MSYNC_1r1w.synth.nz.mem[966] [3];
  assign _05109_ = \bapg_rd.w_ptr_r [1] ? _05108_ : _05107_;
  assign _05110_ = \bapg_rd.w_ptr_r [2] ? _05109_ : _05106_;
  assign _05111_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [3] : \MSYNC_1r1w.synth.nz.mem[968] [3];
  assign _05112_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [3] : \MSYNC_1r1w.synth.nz.mem[970] [3];
  assign _05113_ = \bapg_rd.w_ptr_r [1] ? _05112_ : _05111_;
  assign _05114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [3] : \MSYNC_1r1w.synth.nz.mem[972] [3];
  assign _05115_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [3] : \MSYNC_1r1w.synth.nz.mem[974] [3];
  assign _05116_ = \bapg_rd.w_ptr_r [1] ? _05115_ : _05114_;
  assign _05117_ = \bapg_rd.w_ptr_r [2] ? _05116_ : _05113_;
  assign _05118_ = \bapg_rd.w_ptr_r [3] ? _05117_ : _05110_;
  assign _05119_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [3] : \MSYNC_1r1w.synth.nz.mem[976] [3];
  assign _05120_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [3] : \MSYNC_1r1w.synth.nz.mem[978] [3];
  assign _05121_ = \bapg_rd.w_ptr_r [1] ? _05120_ : _05119_;
  assign _05122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [3] : \MSYNC_1r1w.synth.nz.mem[980] [3];
  assign _05123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [3] : \MSYNC_1r1w.synth.nz.mem[982] [3];
  assign _05124_ = \bapg_rd.w_ptr_r [1] ? _05123_ : _05122_;
  assign _05125_ = \bapg_rd.w_ptr_r [2] ? _05124_ : _05121_;
  assign _05126_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [3] : \MSYNC_1r1w.synth.nz.mem[984] [3];
  assign _05127_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [3] : \MSYNC_1r1w.synth.nz.mem[986] [3];
  assign _05128_ = \bapg_rd.w_ptr_r [1] ? _05127_ : _05126_;
  assign _05129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [3] : \MSYNC_1r1w.synth.nz.mem[988] [3];
  assign _05130_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [3] : \MSYNC_1r1w.synth.nz.mem[990] [3];
  assign _05131_ = \bapg_rd.w_ptr_r [1] ? _05130_ : _05129_;
  assign _05132_ = \bapg_rd.w_ptr_r [2] ? _05131_ : _05128_;
  assign _05133_ = \bapg_rd.w_ptr_r [3] ? _05132_ : _05125_;
  assign _05134_ = \bapg_rd.w_ptr_r [4] ? _05133_ : _05118_;
  assign _05135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [3] : \MSYNC_1r1w.synth.nz.mem[992] [3];
  assign _05136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [3] : \MSYNC_1r1w.synth.nz.mem[994] [3];
  assign _05137_ = \bapg_rd.w_ptr_r [1] ? _05136_ : _05135_;
  assign _05138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [3] : \MSYNC_1r1w.synth.nz.mem[996] [3];
  assign _05139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [3] : \MSYNC_1r1w.synth.nz.mem[998] [3];
  assign _05140_ = \bapg_rd.w_ptr_r [1] ? _05139_ : _05138_;
  assign _05141_ = \bapg_rd.w_ptr_r [2] ? _05140_ : _05137_;
  assign _05142_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [3] : \MSYNC_1r1w.synth.nz.mem[1000] [3];
  assign _05143_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [3] : \MSYNC_1r1w.synth.nz.mem[1002] [3];
  assign _05144_ = \bapg_rd.w_ptr_r [1] ? _05143_ : _05142_;
  assign _05145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [3] : \MSYNC_1r1w.synth.nz.mem[1004] [3];
  assign _05146_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [3] : \MSYNC_1r1w.synth.nz.mem[1006] [3];
  assign _05147_ = \bapg_rd.w_ptr_r [1] ? _05146_ : _05145_;
  assign _05148_ = \bapg_rd.w_ptr_r [2] ? _05147_ : _05144_;
  assign _05149_ = \bapg_rd.w_ptr_r [3] ? _05148_ : _05141_;
  assign _05150_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [3] : \MSYNC_1r1w.synth.nz.mem[1008] [3];
  assign _05151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [3] : \MSYNC_1r1w.synth.nz.mem[1010] [3];
  assign _05152_ = \bapg_rd.w_ptr_r [1] ? _05151_ : _05150_;
  assign _05153_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [3] : \MSYNC_1r1w.synth.nz.mem[1012] [3];
  assign _05154_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [3] : \MSYNC_1r1w.synth.nz.mem[1014] [3];
  assign _05155_ = \bapg_rd.w_ptr_r [1] ? _05154_ : _05153_;
  assign _05156_ = \bapg_rd.w_ptr_r [2] ? _05155_ : _05152_;
  assign _05157_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [3] : \MSYNC_1r1w.synth.nz.mem[1016] [3];
  assign _05158_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [3] : \MSYNC_1r1w.synth.nz.mem[1018] [3];
  assign _05159_ = \bapg_rd.w_ptr_r [1] ? _05158_ : _05157_;
  assign _05160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [3] : \MSYNC_1r1w.synth.nz.mem[1020] [3];
  assign _05161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [3] : \MSYNC_1r1w.synth.nz.mem[1022] [3];
  assign _05162_ = \bapg_rd.w_ptr_r [1] ? _05161_ : _05160_;
  assign _05163_ = \bapg_rd.w_ptr_r [2] ? _05162_ : _05159_;
  assign _05164_ = \bapg_rd.w_ptr_r [3] ? _05163_ : _05156_;
  assign _05165_ = \bapg_rd.w_ptr_r [4] ? _05164_ : _05149_;
  assign _05166_ = \bapg_rd.w_ptr_r [5] ? _05165_ : _05134_;
  assign _05167_ = \bapg_rd.w_ptr_r [6] ? _05166_ : _05103_;
  assign _05168_ = \bapg_rd.w_ptr_r [7] ? _05167_ : _05040_;
  assign _05169_ = \bapg_rd.w_ptr_r [8] ? _05168_ : _04913_;
  assign r_data_o[3] = \bapg_rd.w_ptr_r [9] ? _05169_ : _04658_;
  assign _05170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [4] : \MSYNC_1r1w.synth.nz.mem[0] [4];
  assign _05171_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [4] : \MSYNC_1r1w.synth.nz.mem[2] [4];
  assign _05172_ = \bapg_rd.w_ptr_r [1] ? _05171_ : _05170_;
  assign _05173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [4] : \MSYNC_1r1w.synth.nz.mem[4] [4];
  assign _05174_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [4] : \MSYNC_1r1w.synth.nz.mem[6] [4];
  assign _05175_ = \bapg_rd.w_ptr_r [1] ? _05174_ : _05173_;
  assign _05176_ = \bapg_rd.w_ptr_r [2] ? _05175_ : _05172_;
  assign _05177_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [4] : \MSYNC_1r1w.synth.nz.mem[8] [4];
  assign _05178_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [4] : \MSYNC_1r1w.synth.nz.mem[10] [4];
  assign _05179_ = \bapg_rd.w_ptr_r [1] ? _05178_ : _05177_;
  assign _05180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [4] : \MSYNC_1r1w.synth.nz.mem[12] [4];
  assign _05181_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [4] : \MSYNC_1r1w.synth.nz.mem[14] [4];
  assign _05182_ = \bapg_rd.w_ptr_r [1] ? _05181_ : _05180_;
  assign _05183_ = \bapg_rd.w_ptr_r [2] ? _05182_ : _05179_;
  assign _05184_ = \bapg_rd.w_ptr_r [3] ? _05183_ : _05176_;
  assign _05185_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [4] : \MSYNC_1r1w.synth.nz.mem[16] [4];
  assign _05186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [4] : \MSYNC_1r1w.synth.nz.mem[18] [4];
  assign _05187_ = \bapg_rd.w_ptr_r [1] ? _05186_ : _05185_;
  assign _05188_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [4] : \MSYNC_1r1w.synth.nz.mem[20] [4];
  assign _05189_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [4] : \MSYNC_1r1w.synth.nz.mem[22] [4];
  assign _05190_ = \bapg_rd.w_ptr_r [1] ? _05189_ : _05188_;
  assign _05191_ = \bapg_rd.w_ptr_r [2] ? _05190_ : _05187_;
  assign _05192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [4] : \MSYNC_1r1w.synth.nz.mem[24] [4];
  assign _05193_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [4] : \MSYNC_1r1w.synth.nz.mem[26] [4];
  assign _05194_ = \bapg_rd.w_ptr_r [1] ? _05193_ : _05192_;
  assign _05195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [4] : \MSYNC_1r1w.synth.nz.mem[28] [4];
  assign _05196_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [4] : \MSYNC_1r1w.synth.nz.mem[30] [4];
  assign _05197_ = \bapg_rd.w_ptr_r [1] ? _05196_ : _05195_;
  assign _05198_ = \bapg_rd.w_ptr_r [2] ? _05197_ : _05194_;
  assign _05199_ = \bapg_rd.w_ptr_r [3] ? _05198_ : _05191_;
  assign _05200_ = \bapg_rd.w_ptr_r [4] ? _05199_ : _05184_;
  assign _05201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [4] : \MSYNC_1r1w.synth.nz.mem[32] [4];
  assign _05202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [4] : \MSYNC_1r1w.synth.nz.mem[34] [4];
  assign _05203_ = \bapg_rd.w_ptr_r [1] ? _05202_ : _05201_;
  assign _05204_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [4] : \MSYNC_1r1w.synth.nz.mem[36] [4];
  assign _05205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [4] : \MSYNC_1r1w.synth.nz.mem[38] [4];
  assign _05206_ = \bapg_rd.w_ptr_r [1] ? _05205_ : _05204_;
  assign _05207_ = \bapg_rd.w_ptr_r [2] ? _05206_ : _05203_;
  assign _05208_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [4] : \MSYNC_1r1w.synth.nz.mem[40] [4];
  assign _05209_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [4] : \MSYNC_1r1w.synth.nz.mem[42] [4];
  assign _05210_ = \bapg_rd.w_ptr_r [1] ? _05209_ : _05208_;
  assign _05211_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [4] : \MSYNC_1r1w.synth.nz.mem[44] [4];
  assign _05212_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [4] : \MSYNC_1r1w.synth.nz.mem[46] [4];
  assign _05213_ = \bapg_rd.w_ptr_r [1] ? _05212_ : _05211_;
  assign _05214_ = \bapg_rd.w_ptr_r [2] ? _05213_ : _05210_;
  assign _05215_ = \bapg_rd.w_ptr_r [3] ? _05214_ : _05207_;
  assign _05216_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [4] : \MSYNC_1r1w.synth.nz.mem[48] [4];
  assign _05217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [4] : \MSYNC_1r1w.synth.nz.mem[50] [4];
  assign _05218_ = \bapg_rd.w_ptr_r [1] ? _05217_ : _05216_;
  assign _05219_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [4] : \MSYNC_1r1w.synth.nz.mem[52] [4];
  assign _05220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [4] : \MSYNC_1r1w.synth.nz.mem[54] [4];
  assign _05221_ = \bapg_rd.w_ptr_r [1] ? _05220_ : _05219_;
  assign _05222_ = \bapg_rd.w_ptr_r [2] ? _05221_ : _05218_;
  assign _05223_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [4] : \MSYNC_1r1w.synth.nz.mem[56] [4];
  assign _05224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [4] : \MSYNC_1r1w.synth.nz.mem[58] [4];
  assign _05225_ = \bapg_rd.w_ptr_r [1] ? _05224_ : _05223_;
  assign _05226_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [4] : \MSYNC_1r1w.synth.nz.mem[60] [4];
  assign _05227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [4] : \MSYNC_1r1w.synth.nz.mem[62] [4];
  assign _05228_ = \bapg_rd.w_ptr_r [1] ? _05227_ : _05226_;
  assign _05229_ = \bapg_rd.w_ptr_r [2] ? _05228_ : _05225_;
  assign _05230_ = \bapg_rd.w_ptr_r [3] ? _05229_ : _05222_;
  assign _05231_ = \bapg_rd.w_ptr_r [4] ? _05230_ : _05215_;
  assign _05232_ = \bapg_rd.w_ptr_r [5] ? _05231_ : _05200_;
  assign _05233_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [4] : \MSYNC_1r1w.synth.nz.mem[64] [4];
  assign _05234_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [4] : \MSYNC_1r1w.synth.nz.mem[66] [4];
  assign _05235_ = \bapg_rd.w_ptr_r [1] ? _05234_ : _05233_;
  assign _05236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [4] : \MSYNC_1r1w.synth.nz.mem[68] [4];
  assign _05237_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [4] : \MSYNC_1r1w.synth.nz.mem[70] [4];
  assign _05238_ = \bapg_rd.w_ptr_r [1] ? _05237_ : _05236_;
  assign _05239_ = \bapg_rd.w_ptr_r [2] ? _05238_ : _05235_;
  assign _05240_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [4] : \MSYNC_1r1w.synth.nz.mem[72] [4];
  assign _05241_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [4] : \MSYNC_1r1w.synth.nz.mem[74] [4];
  assign _05242_ = \bapg_rd.w_ptr_r [1] ? _05241_ : _05240_;
  assign _05243_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [4] : \MSYNC_1r1w.synth.nz.mem[76] [4];
  assign _05244_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [4] : \MSYNC_1r1w.synth.nz.mem[78] [4];
  assign _05245_ = \bapg_rd.w_ptr_r [1] ? _05244_ : _05243_;
  assign _05246_ = \bapg_rd.w_ptr_r [2] ? _05245_ : _05242_;
  assign _05247_ = \bapg_rd.w_ptr_r [3] ? _05246_ : _05239_;
  assign _05248_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [4] : \MSYNC_1r1w.synth.nz.mem[80] [4];
  assign _05249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [4] : \MSYNC_1r1w.synth.nz.mem[82] [4];
  assign _05250_ = \bapg_rd.w_ptr_r [1] ? _05249_ : _05248_;
  assign _05251_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [4] : \MSYNC_1r1w.synth.nz.mem[84] [4];
  assign _05252_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [4] : \MSYNC_1r1w.synth.nz.mem[86] [4];
  assign _05253_ = \bapg_rd.w_ptr_r [1] ? _05252_ : _05251_;
  assign _05254_ = \bapg_rd.w_ptr_r [2] ? _05253_ : _05250_;
  assign _05255_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [4] : \MSYNC_1r1w.synth.nz.mem[88] [4];
  assign _05256_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [4] : \MSYNC_1r1w.synth.nz.mem[90] [4];
  assign _05257_ = \bapg_rd.w_ptr_r [1] ? _05256_ : _05255_;
  assign _05258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [4] : \MSYNC_1r1w.synth.nz.mem[92] [4];
  assign _05259_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [4] : \MSYNC_1r1w.synth.nz.mem[94] [4];
  assign _05260_ = \bapg_rd.w_ptr_r [1] ? _05259_ : _05258_;
  assign _05261_ = \bapg_rd.w_ptr_r [2] ? _05260_ : _05257_;
  assign _05262_ = \bapg_rd.w_ptr_r [3] ? _05261_ : _05254_;
  assign _05263_ = \bapg_rd.w_ptr_r [4] ? _05262_ : _05247_;
  assign _05264_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [4] : \MSYNC_1r1w.synth.nz.mem[96] [4];
  assign _05265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [4] : \MSYNC_1r1w.synth.nz.mem[98] [4];
  assign _05266_ = \bapg_rd.w_ptr_r [1] ? _05265_ : _05264_;
  assign _05267_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [4] : \MSYNC_1r1w.synth.nz.mem[100] [4];
  assign _05268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [4] : \MSYNC_1r1w.synth.nz.mem[102] [4];
  assign _05269_ = \bapg_rd.w_ptr_r [1] ? _05268_ : _05267_;
  assign _05270_ = \bapg_rd.w_ptr_r [2] ? _05269_ : _05266_;
  assign _05271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [4] : \MSYNC_1r1w.synth.nz.mem[104] [4];
  assign _05272_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [4] : \MSYNC_1r1w.synth.nz.mem[106] [4];
  assign _05273_ = \bapg_rd.w_ptr_r [1] ? _05272_ : _05271_;
  assign _05274_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [4] : \MSYNC_1r1w.synth.nz.mem[108] [4];
  assign _05275_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [4] : \MSYNC_1r1w.synth.nz.mem[110] [4];
  assign _05276_ = \bapg_rd.w_ptr_r [1] ? _05275_ : _05274_;
  assign _05277_ = \bapg_rd.w_ptr_r [2] ? _05276_ : _05273_;
  assign _05278_ = \bapg_rd.w_ptr_r [3] ? _05277_ : _05270_;
  assign _05279_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [4] : \MSYNC_1r1w.synth.nz.mem[112] [4];
  assign _05280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [4] : \MSYNC_1r1w.synth.nz.mem[114] [4];
  assign _05281_ = \bapg_rd.w_ptr_r [1] ? _05280_ : _05279_;
  assign _05282_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [4] : \MSYNC_1r1w.synth.nz.mem[116] [4];
  assign _05283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [4] : \MSYNC_1r1w.synth.nz.mem[118] [4];
  assign _05284_ = \bapg_rd.w_ptr_r [1] ? _05283_ : _05282_;
  assign _05285_ = \bapg_rd.w_ptr_r [2] ? _05284_ : _05281_;
  assign _05286_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [4] : \MSYNC_1r1w.synth.nz.mem[120] [4];
  assign _05287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [4] : \MSYNC_1r1w.synth.nz.mem[122] [4];
  assign _05288_ = \bapg_rd.w_ptr_r [1] ? _05287_ : _05286_;
  assign _05289_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [4] : \MSYNC_1r1w.synth.nz.mem[124] [4];
  assign _05290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [4] : \MSYNC_1r1w.synth.nz.mem[126] [4];
  assign _05291_ = \bapg_rd.w_ptr_r [1] ? _05290_ : _05289_;
  assign _05292_ = \bapg_rd.w_ptr_r [2] ? _05291_ : _05288_;
  assign _05293_ = \bapg_rd.w_ptr_r [3] ? _05292_ : _05285_;
  assign _05294_ = \bapg_rd.w_ptr_r [4] ? _05293_ : _05278_;
  assign _05295_ = \bapg_rd.w_ptr_r [5] ? _05294_ : _05263_;
  assign _05296_ = \bapg_rd.w_ptr_r [6] ? _05295_ : _05232_;
  assign _05297_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [4] : \MSYNC_1r1w.synth.nz.mem[128] [4];
  assign _05298_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [4] : \MSYNC_1r1w.synth.nz.mem[130] [4];
  assign _05299_ = \bapg_rd.w_ptr_r [1] ? _05298_ : _05297_;
  assign _05300_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [4] : \MSYNC_1r1w.synth.nz.mem[132] [4];
  assign _05301_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [4] : \MSYNC_1r1w.synth.nz.mem[134] [4];
  assign _05302_ = \bapg_rd.w_ptr_r [1] ? _05301_ : _05300_;
  assign _05303_ = \bapg_rd.w_ptr_r [2] ? _05302_ : _05299_;
  assign _05304_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [4] : \MSYNC_1r1w.synth.nz.mem[136] [4];
  assign _05305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [4] : \MSYNC_1r1w.synth.nz.mem[138] [4];
  assign _05306_ = \bapg_rd.w_ptr_r [1] ? _05305_ : _05304_;
  assign _05307_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [4] : \MSYNC_1r1w.synth.nz.mem[140] [4];
  assign _05308_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [4] : \MSYNC_1r1w.synth.nz.mem[142] [4];
  assign _05309_ = \bapg_rd.w_ptr_r [1] ? _05308_ : _05307_;
  assign _05310_ = \bapg_rd.w_ptr_r [2] ? _05309_ : _05306_;
  assign _05311_ = \bapg_rd.w_ptr_r [3] ? _05310_ : _05303_;
  assign _05312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [4] : \MSYNC_1r1w.synth.nz.mem[144] [4];
  assign _05313_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [4] : \MSYNC_1r1w.synth.nz.mem[146] [4];
  assign _05314_ = \bapg_rd.w_ptr_r [1] ? _05313_ : _05312_;
  assign _05315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [4] : \MSYNC_1r1w.synth.nz.mem[148] [4];
  assign _05316_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [4] : \MSYNC_1r1w.synth.nz.mem[150] [4];
  assign _05317_ = \bapg_rd.w_ptr_r [1] ? _05316_ : _05315_;
  assign _05318_ = \bapg_rd.w_ptr_r [2] ? _05317_ : _05314_;
  assign _05319_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [4] : \MSYNC_1r1w.synth.nz.mem[152] [4];
  assign _05320_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [4] : \MSYNC_1r1w.synth.nz.mem[154] [4];
  assign _05321_ = \bapg_rd.w_ptr_r [1] ? _05320_ : _05319_;
  assign _05322_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [4] : \MSYNC_1r1w.synth.nz.mem[156] [4];
  assign _05323_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [4] : \MSYNC_1r1w.synth.nz.mem[158] [4];
  assign _05324_ = \bapg_rd.w_ptr_r [1] ? _05323_ : _05322_;
  assign _05325_ = \bapg_rd.w_ptr_r [2] ? _05324_ : _05321_;
  assign _05326_ = \bapg_rd.w_ptr_r [3] ? _05325_ : _05318_;
  assign _05327_ = \bapg_rd.w_ptr_r [4] ? _05326_ : _05311_;
  assign _05328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [4] : \MSYNC_1r1w.synth.nz.mem[160] [4];
  assign _05329_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [4] : \MSYNC_1r1w.synth.nz.mem[162] [4];
  assign _05330_ = \bapg_rd.w_ptr_r [1] ? _05329_ : _05328_;
  assign _05331_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [4] : \MSYNC_1r1w.synth.nz.mem[164] [4];
  assign _05332_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [4] : \MSYNC_1r1w.synth.nz.mem[166] [4];
  assign _05333_ = \bapg_rd.w_ptr_r [1] ? _05332_ : _05331_;
  assign _05334_ = \bapg_rd.w_ptr_r [2] ? _05333_ : _05330_;
  assign _05335_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [4] : \MSYNC_1r1w.synth.nz.mem[168] [4];
  assign _05336_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [4] : \MSYNC_1r1w.synth.nz.mem[170] [4];
  assign _05337_ = \bapg_rd.w_ptr_r [1] ? _05336_ : _05335_;
  assign _05338_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [4] : \MSYNC_1r1w.synth.nz.mem[172] [4];
  assign _05339_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [4] : \MSYNC_1r1w.synth.nz.mem[174] [4];
  assign _05340_ = \bapg_rd.w_ptr_r [1] ? _05339_ : _05338_;
  assign _05341_ = \bapg_rd.w_ptr_r [2] ? _05340_ : _05337_;
  assign _05342_ = \bapg_rd.w_ptr_r [3] ? _05341_ : _05334_;
  assign _05343_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [4] : \MSYNC_1r1w.synth.nz.mem[176] [4];
  assign _05344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [4] : \MSYNC_1r1w.synth.nz.mem[178] [4];
  assign _05345_ = \bapg_rd.w_ptr_r [1] ? _05344_ : _05343_;
  assign _05346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [4] : \MSYNC_1r1w.synth.nz.mem[180] [4];
  assign _05347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [4] : \MSYNC_1r1w.synth.nz.mem[182] [4];
  assign _05348_ = \bapg_rd.w_ptr_r [1] ? _05347_ : _05346_;
  assign _05349_ = \bapg_rd.w_ptr_r [2] ? _05348_ : _05345_;
  assign _05350_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [4] : \MSYNC_1r1w.synth.nz.mem[184] [4];
  assign _05351_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [4] : \MSYNC_1r1w.synth.nz.mem[186] [4];
  assign _05352_ = \bapg_rd.w_ptr_r [1] ? _05351_ : _05350_;
  assign _05353_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [4] : \MSYNC_1r1w.synth.nz.mem[188] [4];
  assign _05354_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [4] : \MSYNC_1r1w.synth.nz.mem[190] [4];
  assign _05355_ = \bapg_rd.w_ptr_r [1] ? _05354_ : _05353_;
  assign _05356_ = \bapg_rd.w_ptr_r [2] ? _05355_ : _05352_;
  assign _05357_ = \bapg_rd.w_ptr_r [3] ? _05356_ : _05349_;
  assign _05358_ = \bapg_rd.w_ptr_r [4] ? _05357_ : _05342_;
  assign _05359_ = \bapg_rd.w_ptr_r [5] ? _05358_ : _05327_;
  assign _05360_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [4] : \MSYNC_1r1w.synth.nz.mem[192] [4];
  assign _05361_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [4] : \MSYNC_1r1w.synth.nz.mem[194] [4];
  assign _05362_ = \bapg_rd.w_ptr_r [1] ? _05361_ : _05360_;
  assign _05363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [4] : \MSYNC_1r1w.synth.nz.mem[196] [4];
  assign _05364_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [4] : \MSYNC_1r1w.synth.nz.mem[198] [4];
  assign _05365_ = \bapg_rd.w_ptr_r [1] ? _05364_ : _05363_;
  assign _05366_ = \bapg_rd.w_ptr_r [2] ? _05365_ : _05362_;
  assign _05367_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [4] : \MSYNC_1r1w.synth.nz.mem[200] [4];
  assign _05368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [4] : \MSYNC_1r1w.synth.nz.mem[202] [4];
  assign _05369_ = \bapg_rd.w_ptr_r [1] ? _05368_ : _05367_;
  assign _05370_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [4] : \MSYNC_1r1w.synth.nz.mem[204] [4];
  assign _05371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [4] : \MSYNC_1r1w.synth.nz.mem[206] [4];
  assign _05372_ = \bapg_rd.w_ptr_r [1] ? _05371_ : _05370_;
  assign _05373_ = \bapg_rd.w_ptr_r [2] ? _05372_ : _05369_;
  assign _05374_ = \bapg_rd.w_ptr_r [3] ? _05373_ : _05366_;
  assign _05375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [4] : \MSYNC_1r1w.synth.nz.mem[208] [4];
  assign _05376_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [4] : \MSYNC_1r1w.synth.nz.mem[210] [4];
  assign _05377_ = \bapg_rd.w_ptr_r [1] ? _05376_ : _05375_;
  assign _05378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [4] : \MSYNC_1r1w.synth.nz.mem[212] [4];
  assign _05379_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [4] : \MSYNC_1r1w.synth.nz.mem[214] [4];
  assign _05380_ = \bapg_rd.w_ptr_r [1] ? _05379_ : _05378_;
  assign _05381_ = \bapg_rd.w_ptr_r [2] ? _05380_ : _05377_;
  assign _05382_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [4] : \MSYNC_1r1w.synth.nz.mem[216] [4];
  assign _05383_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [4] : \MSYNC_1r1w.synth.nz.mem[218] [4];
  assign _05384_ = \bapg_rd.w_ptr_r [1] ? _05383_ : _05382_;
  assign _05385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [4] : \MSYNC_1r1w.synth.nz.mem[220] [4];
  assign _05386_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [4] : \MSYNC_1r1w.synth.nz.mem[222] [4];
  assign _05387_ = \bapg_rd.w_ptr_r [1] ? _05386_ : _05385_;
  assign _05388_ = \bapg_rd.w_ptr_r [2] ? _05387_ : _05384_;
  assign _05389_ = \bapg_rd.w_ptr_r [3] ? _05388_ : _05381_;
  assign _05390_ = \bapg_rd.w_ptr_r [4] ? _05389_ : _05374_;
  assign _05391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [4] : \MSYNC_1r1w.synth.nz.mem[224] [4];
  assign _05392_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [4] : \MSYNC_1r1w.synth.nz.mem[226] [4];
  assign _05393_ = \bapg_rd.w_ptr_r [1] ? _05392_ : _05391_;
  assign _05394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [4] : \MSYNC_1r1w.synth.nz.mem[228] [4];
  assign _05395_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [4] : \MSYNC_1r1w.synth.nz.mem[230] [4];
  assign _05396_ = \bapg_rd.w_ptr_r [1] ? _05395_ : _05394_;
  assign _05397_ = \bapg_rd.w_ptr_r [2] ? _05396_ : _05393_;
  assign _05398_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [4] : \MSYNC_1r1w.synth.nz.mem[232] [4];
  assign _05399_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [4] : \MSYNC_1r1w.synth.nz.mem[234] [4];
  assign _05400_ = \bapg_rd.w_ptr_r [1] ? _05399_ : _05398_;
  assign _05401_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [4] : \MSYNC_1r1w.synth.nz.mem[236] [4];
  assign _05402_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [4] : \MSYNC_1r1w.synth.nz.mem[238] [4];
  assign _05403_ = \bapg_rd.w_ptr_r [1] ? _05402_ : _05401_;
  assign _05404_ = \bapg_rd.w_ptr_r [2] ? _05403_ : _05400_;
  assign _05405_ = \bapg_rd.w_ptr_r [3] ? _05404_ : _05397_;
  assign _05406_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [4] : \MSYNC_1r1w.synth.nz.mem[240] [4];
  assign _05407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [4] : \MSYNC_1r1w.synth.nz.mem[242] [4];
  assign _05408_ = \bapg_rd.w_ptr_r [1] ? _05407_ : _05406_;
  assign _05409_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [4] : \MSYNC_1r1w.synth.nz.mem[244] [4];
  assign _05410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [4] : \MSYNC_1r1w.synth.nz.mem[246] [4];
  assign _05411_ = \bapg_rd.w_ptr_r [1] ? _05410_ : _05409_;
  assign _05412_ = \bapg_rd.w_ptr_r [2] ? _05411_ : _05408_;
  assign _05413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [4] : \MSYNC_1r1w.synth.nz.mem[248] [4];
  assign _05414_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [4] : \MSYNC_1r1w.synth.nz.mem[250] [4];
  assign _05415_ = \bapg_rd.w_ptr_r [1] ? _05414_ : _05413_;
  assign _05416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [4] : \MSYNC_1r1w.synth.nz.mem[252] [4];
  assign _05417_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [4] : \MSYNC_1r1w.synth.nz.mem[254] [4];
  assign _05418_ = \bapg_rd.w_ptr_r [1] ? _05417_ : _05416_;
  assign _05419_ = \bapg_rd.w_ptr_r [2] ? _05418_ : _05415_;
  assign _05420_ = \bapg_rd.w_ptr_r [3] ? _05419_ : _05412_;
  assign _05421_ = \bapg_rd.w_ptr_r [4] ? _05420_ : _05405_;
  assign _05422_ = \bapg_rd.w_ptr_r [5] ? _05421_ : _05390_;
  assign _05423_ = \bapg_rd.w_ptr_r [6] ? _05422_ : _05359_;
  assign _05424_ = \bapg_rd.w_ptr_r [7] ? _05423_ : _05296_;
  assign _05425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [4] : \MSYNC_1r1w.synth.nz.mem[256] [4];
  assign _05426_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [4] : \MSYNC_1r1w.synth.nz.mem[258] [4];
  assign _05427_ = \bapg_rd.w_ptr_r [1] ? _05426_ : _05425_;
  assign _05428_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [4] : \MSYNC_1r1w.synth.nz.mem[260] [4];
  assign _05429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [4] : \MSYNC_1r1w.synth.nz.mem[262] [4];
  assign _05430_ = \bapg_rd.w_ptr_r [1] ? _05429_ : _05428_;
  assign _05431_ = \bapg_rd.w_ptr_r [2] ? _05430_ : _05427_;
  assign _05432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [4] : \MSYNC_1r1w.synth.nz.mem[264] [4];
  assign _05433_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [4] : \MSYNC_1r1w.synth.nz.mem[266] [4];
  assign _05434_ = \bapg_rd.w_ptr_r [1] ? _05433_ : _05432_;
  assign _05435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [4] : \MSYNC_1r1w.synth.nz.mem[268] [4];
  assign _05436_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [4] : \MSYNC_1r1w.synth.nz.mem[270] [4];
  assign _05437_ = \bapg_rd.w_ptr_r [1] ? _05436_ : _05435_;
  assign _05438_ = \bapg_rd.w_ptr_r [2] ? _05437_ : _05434_;
  assign _05439_ = \bapg_rd.w_ptr_r [3] ? _05438_ : _05431_;
  assign _05440_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [4] : \MSYNC_1r1w.synth.nz.mem[272] [4];
  assign _05441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [4] : \MSYNC_1r1w.synth.nz.mem[274] [4];
  assign _05442_ = \bapg_rd.w_ptr_r [1] ? _05441_ : _05440_;
  assign _05443_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [4] : \MSYNC_1r1w.synth.nz.mem[276] [4];
  assign _05444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [4] : \MSYNC_1r1w.synth.nz.mem[278] [4];
  assign _05445_ = \bapg_rd.w_ptr_r [1] ? _05444_ : _05443_;
  assign _05446_ = \bapg_rd.w_ptr_r [2] ? _05445_ : _05442_;
  assign _05447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [4] : \MSYNC_1r1w.synth.nz.mem[280] [4];
  assign _05448_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [4] : \MSYNC_1r1w.synth.nz.mem[282] [4];
  assign _05449_ = \bapg_rd.w_ptr_r [1] ? _05448_ : _05447_;
  assign _05450_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [4] : \MSYNC_1r1w.synth.nz.mem[284] [4];
  assign _05451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [4] : \MSYNC_1r1w.synth.nz.mem[286] [4];
  assign _05452_ = \bapg_rd.w_ptr_r [1] ? _05451_ : _05450_;
  assign _05453_ = \bapg_rd.w_ptr_r [2] ? _05452_ : _05449_;
  assign _05454_ = \bapg_rd.w_ptr_r [3] ? _05453_ : _05446_;
  assign _05455_ = \bapg_rd.w_ptr_r [4] ? _05454_ : _05439_;
  assign _05456_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [4] : \MSYNC_1r1w.synth.nz.mem[288] [4];
  assign _05457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [4] : \MSYNC_1r1w.synth.nz.mem[290] [4];
  assign _05458_ = \bapg_rd.w_ptr_r [1] ? _05457_ : _05456_;
  assign _05459_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [4] : \MSYNC_1r1w.synth.nz.mem[292] [4];
  assign _05460_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [4] : \MSYNC_1r1w.synth.nz.mem[294] [4];
  assign _05461_ = \bapg_rd.w_ptr_r [1] ? _05460_ : _05459_;
  assign _05462_ = \bapg_rd.w_ptr_r [2] ? _05461_ : _05458_;
  assign _05463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [4] : \MSYNC_1r1w.synth.nz.mem[296] [4];
  assign _05464_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [4] : \MSYNC_1r1w.synth.nz.mem[298] [4];
  assign _05465_ = \bapg_rd.w_ptr_r [1] ? _05464_ : _05463_;
  assign _05466_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [4] : \MSYNC_1r1w.synth.nz.mem[300] [4];
  assign _05467_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [4] : \MSYNC_1r1w.synth.nz.mem[302] [4];
  assign _05468_ = \bapg_rd.w_ptr_r [1] ? _05467_ : _05466_;
  assign _05469_ = \bapg_rd.w_ptr_r [2] ? _05468_ : _05465_;
  assign _05470_ = \bapg_rd.w_ptr_r [3] ? _05469_ : _05462_;
  assign _05471_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [4] : \MSYNC_1r1w.synth.nz.mem[304] [4];
  assign _05472_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [4] : \MSYNC_1r1w.synth.nz.mem[306] [4];
  assign _05473_ = \bapg_rd.w_ptr_r [1] ? _05472_ : _05471_;
  assign _05474_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [4] : \MSYNC_1r1w.synth.nz.mem[308] [4];
  assign _05475_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [4] : \MSYNC_1r1w.synth.nz.mem[310] [4];
  assign _05476_ = \bapg_rd.w_ptr_r [1] ? _05475_ : _05474_;
  assign _05477_ = \bapg_rd.w_ptr_r [2] ? _05476_ : _05473_;
  assign _05478_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [4] : \MSYNC_1r1w.synth.nz.mem[312] [4];
  assign _05479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [4] : \MSYNC_1r1w.synth.nz.mem[314] [4];
  assign _05480_ = \bapg_rd.w_ptr_r [1] ? _05479_ : _05478_;
  assign _05481_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [4] : \MSYNC_1r1w.synth.nz.mem[316] [4];
  assign _05482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [4] : \MSYNC_1r1w.synth.nz.mem[318] [4];
  assign _05483_ = \bapg_rd.w_ptr_r [1] ? _05482_ : _05481_;
  assign _05484_ = \bapg_rd.w_ptr_r [2] ? _05483_ : _05480_;
  assign _05485_ = \bapg_rd.w_ptr_r [3] ? _05484_ : _05477_;
  assign _05486_ = \bapg_rd.w_ptr_r [4] ? _05485_ : _05470_;
  assign _05487_ = \bapg_rd.w_ptr_r [5] ? _05486_ : _05455_;
  assign _05488_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [4] : \MSYNC_1r1w.synth.nz.mem[320] [4];
  assign _05489_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [4] : \MSYNC_1r1w.synth.nz.mem[322] [4];
  assign _05490_ = \bapg_rd.w_ptr_r [1] ? _05489_ : _05488_;
  assign _05491_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [4] : \MSYNC_1r1w.synth.nz.mem[324] [4];
  assign _05492_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [4] : \MSYNC_1r1w.synth.nz.mem[326] [4];
  assign _05493_ = \bapg_rd.w_ptr_r [1] ? _05492_ : _05491_;
  assign _05494_ = \bapg_rd.w_ptr_r [2] ? _05493_ : _05490_;
  assign _05495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [4] : \MSYNC_1r1w.synth.nz.mem[328] [4];
  assign _05496_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [4] : \MSYNC_1r1w.synth.nz.mem[330] [4];
  assign _05497_ = \bapg_rd.w_ptr_r [1] ? _05496_ : _05495_;
  assign _05498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [4] : \MSYNC_1r1w.synth.nz.mem[332] [4];
  assign _05499_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [4] : \MSYNC_1r1w.synth.nz.mem[334] [4];
  assign _05500_ = \bapg_rd.w_ptr_r [1] ? _05499_ : _05498_;
  assign _05501_ = \bapg_rd.w_ptr_r [2] ? _05500_ : _05497_;
  assign _05502_ = \bapg_rd.w_ptr_r [3] ? _05501_ : _05494_;
  assign _05503_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [4] : \MSYNC_1r1w.synth.nz.mem[336] [4];
  assign _05504_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [4] : \MSYNC_1r1w.synth.nz.mem[338] [4];
  assign _05505_ = \bapg_rd.w_ptr_r [1] ? _05504_ : _05503_;
  assign _05506_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [4] : \MSYNC_1r1w.synth.nz.mem[340] [4];
  assign _05507_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [4] : \MSYNC_1r1w.synth.nz.mem[342] [4];
  assign _05508_ = \bapg_rd.w_ptr_r [1] ? _05507_ : _05506_;
  assign _05509_ = \bapg_rd.w_ptr_r [2] ? _05508_ : _05505_;
  assign _05510_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [4] : \MSYNC_1r1w.synth.nz.mem[344] [4];
  assign _05511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [4] : \MSYNC_1r1w.synth.nz.mem[346] [4];
  assign _05512_ = \bapg_rd.w_ptr_r [1] ? _05511_ : _05510_;
  assign _05513_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [4] : \MSYNC_1r1w.synth.nz.mem[348] [4];
  assign _05514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [4] : \MSYNC_1r1w.synth.nz.mem[350] [4];
  assign _05515_ = \bapg_rd.w_ptr_r [1] ? _05514_ : _05513_;
  assign _05516_ = \bapg_rd.w_ptr_r [2] ? _05515_ : _05512_;
  assign _05517_ = \bapg_rd.w_ptr_r [3] ? _05516_ : _05509_;
  assign _05518_ = \bapg_rd.w_ptr_r [4] ? _05517_ : _05502_;
  assign _05519_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [4] : \MSYNC_1r1w.synth.nz.mem[352] [4];
  assign _05520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [4] : \MSYNC_1r1w.synth.nz.mem[354] [4];
  assign _05521_ = \bapg_rd.w_ptr_r [1] ? _05520_ : _05519_;
  assign _05522_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [4] : \MSYNC_1r1w.synth.nz.mem[356] [4];
  assign _05523_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [4] : \MSYNC_1r1w.synth.nz.mem[358] [4];
  assign _05524_ = \bapg_rd.w_ptr_r [1] ? _05523_ : _05522_;
  assign _05525_ = \bapg_rd.w_ptr_r [2] ? _05524_ : _05521_;
  assign _05526_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [4] : \MSYNC_1r1w.synth.nz.mem[360] [4];
  assign _05527_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [4] : \MSYNC_1r1w.synth.nz.mem[362] [4];
  assign _05528_ = \bapg_rd.w_ptr_r [1] ? _05527_ : _05526_;
  assign _05529_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [4] : \MSYNC_1r1w.synth.nz.mem[364] [4];
  assign _05530_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [4] : \MSYNC_1r1w.synth.nz.mem[366] [4];
  assign _05531_ = \bapg_rd.w_ptr_r [1] ? _05530_ : _05529_;
  assign _05532_ = \bapg_rd.w_ptr_r [2] ? _05531_ : _05528_;
  assign _05533_ = \bapg_rd.w_ptr_r [3] ? _05532_ : _05525_;
  assign _05534_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [4] : \MSYNC_1r1w.synth.nz.mem[368] [4];
  assign _05535_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [4] : \MSYNC_1r1w.synth.nz.mem[370] [4];
  assign _05536_ = \bapg_rd.w_ptr_r [1] ? _05535_ : _05534_;
  assign _05537_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [4] : \MSYNC_1r1w.synth.nz.mem[372] [4];
  assign _05538_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [4] : \MSYNC_1r1w.synth.nz.mem[374] [4];
  assign _05539_ = \bapg_rd.w_ptr_r [1] ? _05538_ : _05537_;
  assign _05540_ = \bapg_rd.w_ptr_r [2] ? _05539_ : _05536_;
  assign _05541_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [4] : \MSYNC_1r1w.synth.nz.mem[376] [4];
  assign _05542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [4] : \MSYNC_1r1w.synth.nz.mem[378] [4];
  assign _05543_ = \bapg_rd.w_ptr_r [1] ? _05542_ : _05541_;
  assign _05544_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [4] : \MSYNC_1r1w.synth.nz.mem[380] [4];
  assign _05545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [4] : \MSYNC_1r1w.synth.nz.mem[382] [4];
  assign _05546_ = \bapg_rd.w_ptr_r [1] ? _05545_ : _05544_;
  assign _05547_ = \bapg_rd.w_ptr_r [2] ? _05546_ : _05543_;
  assign _05548_ = \bapg_rd.w_ptr_r [3] ? _05547_ : _05540_;
  assign _05549_ = \bapg_rd.w_ptr_r [4] ? _05548_ : _05533_;
  assign _05550_ = \bapg_rd.w_ptr_r [5] ? _05549_ : _05518_;
  assign _05551_ = \bapg_rd.w_ptr_r [6] ? _05550_ : _05487_;
  assign _05552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [4] : \MSYNC_1r1w.synth.nz.mem[384] [4];
  assign _05553_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [4] : \MSYNC_1r1w.synth.nz.mem[386] [4];
  assign _05554_ = \bapg_rd.w_ptr_r [1] ? _05553_ : _05552_;
  assign _05555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [4] : \MSYNC_1r1w.synth.nz.mem[388] [4];
  assign _05556_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [4] : \MSYNC_1r1w.synth.nz.mem[390] [4];
  assign _05557_ = \bapg_rd.w_ptr_r [1] ? _05556_ : _05555_;
  assign _05558_ = \bapg_rd.w_ptr_r [2] ? _05557_ : _05554_;
  assign _05559_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [4] : \MSYNC_1r1w.synth.nz.mem[392] [4];
  assign _05560_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [4] : \MSYNC_1r1w.synth.nz.mem[394] [4];
  assign _05561_ = \bapg_rd.w_ptr_r [1] ? _05560_ : _05559_;
  assign _05562_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [4] : \MSYNC_1r1w.synth.nz.mem[396] [4];
  assign _05563_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [4] : \MSYNC_1r1w.synth.nz.mem[398] [4];
  assign _05564_ = \bapg_rd.w_ptr_r [1] ? _05563_ : _05562_;
  assign _05565_ = \bapg_rd.w_ptr_r [2] ? _05564_ : _05561_;
  assign _05566_ = \bapg_rd.w_ptr_r [3] ? _05565_ : _05558_;
  assign _05567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [4] : \MSYNC_1r1w.synth.nz.mem[400] [4];
  assign _05568_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [4] : \MSYNC_1r1w.synth.nz.mem[402] [4];
  assign _05569_ = \bapg_rd.w_ptr_r [1] ? _05568_ : _05567_;
  assign _05570_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [4] : \MSYNC_1r1w.synth.nz.mem[404] [4];
  assign _05571_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [4] : \MSYNC_1r1w.synth.nz.mem[406] [4];
  assign _05572_ = \bapg_rd.w_ptr_r [1] ? _05571_ : _05570_;
  assign _05573_ = \bapg_rd.w_ptr_r [2] ? _05572_ : _05569_;
  assign _05574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [4] : \MSYNC_1r1w.synth.nz.mem[408] [4];
  assign _05575_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [4] : \MSYNC_1r1w.synth.nz.mem[410] [4];
  assign _05576_ = \bapg_rd.w_ptr_r [1] ? _05575_ : _05574_;
  assign _05577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [4] : \MSYNC_1r1w.synth.nz.mem[412] [4];
  assign _05578_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [4] : \MSYNC_1r1w.synth.nz.mem[414] [4];
  assign _05579_ = \bapg_rd.w_ptr_r [1] ? _05578_ : _05577_;
  assign _05580_ = \bapg_rd.w_ptr_r [2] ? _05579_ : _05576_;
  assign _05581_ = \bapg_rd.w_ptr_r [3] ? _05580_ : _05573_;
  assign _05582_ = \bapg_rd.w_ptr_r [4] ? _05581_ : _05566_;
  assign _05583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [4] : \MSYNC_1r1w.synth.nz.mem[416] [4];
  assign _05584_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [4] : \MSYNC_1r1w.synth.nz.mem[418] [4];
  assign _05585_ = \bapg_rd.w_ptr_r [1] ? _05584_ : _05583_;
  assign _05586_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [4] : \MSYNC_1r1w.synth.nz.mem[420] [4];
  assign _05587_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [4] : \MSYNC_1r1w.synth.nz.mem[422] [4];
  assign _05588_ = \bapg_rd.w_ptr_r [1] ? _05587_ : _05586_;
  assign _05589_ = \bapg_rd.w_ptr_r [2] ? _05588_ : _05585_;
  assign _05590_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [4] : \MSYNC_1r1w.synth.nz.mem[424] [4];
  assign _05591_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [4] : \MSYNC_1r1w.synth.nz.mem[426] [4];
  assign _05592_ = \bapg_rd.w_ptr_r [1] ? _05591_ : _05590_;
  assign _05593_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [4] : \MSYNC_1r1w.synth.nz.mem[428] [4];
  assign _05594_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [4] : \MSYNC_1r1w.synth.nz.mem[430] [4];
  assign _05595_ = \bapg_rd.w_ptr_r [1] ? _05594_ : _05593_;
  assign _05596_ = \bapg_rd.w_ptr_r [2] ? _05595_ : _05592_;
  assign _05597_ = \bapg_rd.w_ptr_r [3] ? _05596_ : _05589_;
  assign _05598_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [4] : \MSYNC_1r1w.synth.nz.mem[432] [4];
  assign _05599_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [4] : \MSYNC_1r1w.synth.nz.mem[434] [4];
  assign _05600_ = \bapg_rd.w_ptr_r [1] ? _05599_ : _05598_;
  assign _05601_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [4] : \MSYNC_1r1w.synth.nz.mem[436] [4];
  assign _05602_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [4] : \MSYNC_1r1w.synth.nz.mem[438] [4];
  assign _05603_ = \bapg_rd.w_ptr_r [1] ? _05602_ : _05601_;
  assign _05604_ = \bapg_rd.w_ptr_r [2] ? _05603_ : _05600_;
  assign _05605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [4] : \MSYNC_1r1w.synth.nz.mem[440] [4];
  assign _05606_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [4] : \MSYNC_1r1w.synth.nz.mem[442] [4];
  assign _05607_ = \bapg_rd.w_ptr_r [1] ? _05606_ : _05605_;
  assign _05608_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [4] : \MSYNC_1r1w.synth.nz.mem[444] [4];
  assign _05609_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [4] : \MSYNC_1r1w.synth.nz.mem[446] [4];
  assign _05610_ = \bapg_rd.w_ptr_r [1] ? _05609_ : _05608_;
  assign _05611_ = \bapg_rd.w_ptr_r [2] ? _05610_ : _05607_;
  assign _05612_ = \bapg_rd.w_ptr_r [3] ? _05611_ : _05604_;
  assign _05613_ = \bapg_rd.w_ptr_r [4] ? _05612_ : _05597_;
  assign _05614_ = \bapg_rd.w_ptr_r [5] ? _05613_ : _05582_;
  assign _05615_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [4] : \MSYNC_1r1w.synth.nz.mem[448] [4];
  assign _05616_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [4] : \MSYNC_1r1w.synth.nz.mem[450] [4];
  assign _05617_ = \bapg_rd.w_ptr_r [1] ? _05616_ : _05615_;
  assign _05618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [4] : \MSYNC_1r1w.synth.nz.mem[452] [4];
  assign _05619_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [4] : \MSYNC_1r1w.synth.nz.mem[454] [4];
  assign _05620_ = \bapg_rd.w_ptr_r [1] ? _05619_ : _05618_;
  assign _05621_ = \bapg_rd.w_ptr_r [2] ? _05620_ : _05617_;
  assign _05622_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [4] : \MSYNC_1r1w.synth.nz.mem[456] [4];
  assign _05623_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [4] : \MSYNC_1r1w.synth.nz.mem[458] [4];
  assign _05624_ = \bapg_rd.w_ptr_r [1] ? _05623_ : _05622_;
  assign _05625_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [4] : \MSYNC_1r1w.synth.nz.mem[460] [4];
  assign _05626_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [4] : \MSYNC_1r1w.synth.nz.mem[462] [4];
  assign _05627_ = \bapg_rd.w_ptr_r [1] ? _05626_ : _05625_;
  assign _05628_ = \bapg_rd.w_ptr_r [2] ? _05627_ : _05624_;
  assign _05629_ = \bapg_rd.w_ptr_r [3] ? _05628_ : _05621_;
  assign _05630_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [4] : \MSYNC_1r1w.synth.nz.mem[464] [4];
  assign _05631_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [4] : \MSYNC_1r1w.synth.nz.mem[466] [4];
  assign _05632_ = \bapg_rd.w_ptr_r [1] ? _05631_ : _05630_;
  assign _05633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [4] : \MSYNC_1r1w.synth.nz.mem[468] [4];
  assign _05634_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [4] : \MSYNC_1r1w.synth.nz.mem[470] [4];
  assign _05635_ = \bapg_rd.w_ptr_r [1] ? _05634_ : _05633_;
  assign _05636_ = \bapg_rd.w_ptr_r [2] ? _05635_ : _05632_;
  assign _05637_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [4] : \MSYNC_1r1w.synth.nz.mem[472] [4];
  assign _05638_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [4] : \MSYNC_1r1w.synth.nz.mem[474] [4];
  assign _05639_ = \bapg_rd.w_ptr_r [1] ? _05638_ : _05637_;
  assign _05640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [4] : \MSYNC_1r1w.synth.nz.mem[476] [4];
  assign _05641_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [4] : \MSYNC_1r1w.synth.nz.mem[478] [4];
  assign _05642_ = \bapg_rd.w_ptr_r [1] ? _05641_ : _05640_;
  assign _05643_ = \bapg_rd.w_ptr_r [2] ? _05642_ : _05639_;
  assign _05644_ = \bapg_rd.w_ptr_r [3] ? _05643_ : _05636_;
  assign _05645_ = \bapg_rd.w_ptr_r [4] ? _05644_ : _05629_;
  assign _05646_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [4] : \MSYNC_1r1w.synth.nz.mem[480] [4];
  assign _05647_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [4] : \MSYNC_1r1w.synth.nz.mem[482] [4];
  assign _05648_ = \bapg_rd.w_ptr_r [1] ? _05647_ : _05646_;
  assign _05649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [4] : \MSYNC_1r1w.synth.nz.mem[484] [4];
  assign _05650_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [4] : \MSYNC_1r1w.synth.nz.mem[486] [4];
  assign _05651_ = \bapg_rd.w_ptr_r [1] ? _05650_ : _05649_;
  assign _05652_ = \bapg_rd.w_ptr_r [2] ? _05651_ : _05648_;
  assign _05653_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [4] : \MSYNC_1r1w.synth.nz.mem[488] [4];
  assign _05654_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [4] : \MSYNC_1r1w.synth.nz.mem[490] [4];
  assign _05655_ = \bapg_rd.w_ptr_r [1] ? _05654_ : _05653_;
  assign _05656_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [4] : \MSYNC_1r1w.synth.nz.mem[492] [4];
  assign _05657_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [4] : \MSYNC_1r1w.synth.nz.mem[494] [4];
  assign _05658_ = \bapg_rd.w_ptr_r [1] ? _05657_ : _05656_;
  assign _05659_ = \bapg_rd.w_ptr_r [2] ? _05658_ : _05655_;
  assign _05660_ = \bapg_rd.w_ptr_r [3] ? _05659_ : _05652_;
  assign _05661_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [4] : \MSYNC_1r1w.synth.nz.mem[496] [4];
  assign _05662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [4] : \MSYNC_1r1w.synth.nz.mem[498] [4];
  assign _05663_ = \bapg_rd.w_ptr_r [1] ? _05662_ : _05661_;
  assign _05664_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [4] : \MSYNC_1r1w.synth.nz.mem[500] [4];
  assign _05665_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [4] : \MSYNC_1r1w.synth.nz.mem[502] [4];
  assign _05666_ = \bapg_rd.w_ptr_r [1] ? _05665_ : _05664_;
  assign _05667_ = \bapg_rd.w_ptr_r [2] ? _05666_ : _05663_;
  assign _05668_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [4] : \MSYNC_1r1w.synth.nz.mem[504] [4];
  assign _05669_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [4] : \MSYNC_1r1w.synth.nz.mem[506] [4];
  assign _05670_ = \bapg_rd.w_ptr_r [1] ? _05669_ : _05668_;
  assign _05671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [4] : \MSYNC_1r1w.synth.nz.mem[508] [4];
  assign _05672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [4] : \MSYNC_1r1w.synth.nz.mem[510] [4];
  assign _05673_ = \bapg_rd.w_ptr_r [1] ? _05672_ : _05671_;
  assign _05674_ = \bapg_rd.w_ptr_r [2] ? _05673_ : _05670_;
  assign _05675_ = \bapg_rd.w_ptr_r [3] ? _05674_ : _05667_;
  assign _05676_ = \bapg_rd.w_ptr_r [4] ? _05675_ : _05660_;
  assign _05677_ = \bapg_rd.w_ptr_r [5] ? _05676_ : _05645_;
  assign _05678_ = \bapg_rd.w_ptr_r [6] ? _05677_ : _05614_;
  assign _05679_ = \bapg_rd.w_ptr_r [7] ? _05678_ : _05551_;
  assign _05680_ = \bapg_rd.w_ptr_r [8] ? _05679_ : _05424_;
  assign _05681_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [4] : \MSYNC_1r1w.synth.nz.mem[512] [4];
  assign _05682_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [4] : \MSYNC_1r1w.synth.nz.mem[514] [4];
  assign _05683_ = \bapg_rd.w_ptr_r [1] ? _05682_ : _05681_;
  assign _05684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [4] : \MSYNC_1r1w.synth.nz.mem[516] [4];
  assign _05685_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [4] : \MSYNC_1r1w.synth.nz.mem[518] [4];
  assign _05686_ = \bapg_rd.w_ptr_r [1] ? _05685_ : _05684_;
  assign _05687_ = \bapg_rd.w_ptr_r [2] ? _05686_ : _05683_;
  assign _05688_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [4] : \MSYNC_1r1w.synth.nz.mem[520] [4];
  assign _05689_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [4] : \MSYNC_1r1w.synth.nz.mem[522] [4];
  assign _05690_ = \bapg_rd.w_ptr_r [1] ? _05689_ : _05688_;
  assign _05691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [4] : \MSYNC_1r1w.synth.nz.mem[524] [4];
  assign _05692_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [4] : \MSYNC_1r1w.synth.nz.mem[526] [4];
  assign _05693_ = \bapg_rd.w_ptr_r [1] ? _05692_ : _05691_;
  assign _05694_ = \bapg_rd.w_ptr_r [2] ? _05693_ : _05690_;
  assign _05695_ = \bapg_rd.w_ptr_r [3] ? _05694_ : _05687_;
  assign _05696_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [4] : \MSYNC_1r1w.synth.nz.mem[528] [4];
  assign _05697_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [4] : \MSYNC_1r1w.synth.nz.mem[530] [4];
  assign _05698_ = \bapg_rd.w_ptr_r [1] ? _05697_ : _05696_;
  assign _05699_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [4] : \MSYNC_1r1w.synth.nz.mem[532] [4];
  assign _05700_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [4] : \MSYNC_1r1w.synth.nz.mem[534] [4];
  assign _05701_ = \bapg_rd.w_ptr_r [1] ? _05700_ : _05699_;
  assign _05702_ = \bapg_rd.w_ptr_r [2] ? _05701_ : _05698_;
  assign _05703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [4] : \MSYNC_1r1w.synth.nz.mem[536] [4];
  assign _05704_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [4] : \MSYNC_1r1w.synth.nz.mem[538] [4];
  assign _05705_ = \bapg_rd.w_ptr_r [1] ? _05704_ : _05703_;
  assign _05706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [4] : \MSYNC_1r1w.synth.nz.mem[540] [4];
  assign _05707_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [4] : \MSYNC_1r1w.synth.nz.mem[542] [4];
  assign _05708_ = \bapg_rd.w_ptr_r [1] ? _05707_ : _05706_;
  assign _05709_ = \bapg_rd.w_ptr_r [2] ? _05708_ : _05705_;
  assign _05710_ = \bapg_rd.w_ptr_r [3] ? _05709_ : _05702_;
  assign _05711_ = \bapg_rd.w_ptr_r [4] ? _05710_ : _05695_;
  assign _05712_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [4] : \MSYNC_1r1w.synth.nz.mem[544] [4];
  assign _05713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [4] : \MSYNC_1r1w.synth.nz.mem[546] [4];
  assign _05714_ = \bapg_rd.w_ptr_r [1] ? _05713_ : _05712_;
  assign _05715_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [4] : \MSYNC_1r1w.synth.nz.mem[548] [4];
  assign _05716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [4] : \MSYNC_1r1w.synth.nz.mem[550] [4];
  assign _05717_ = \bapg_rd.w_ptr_r [1] ? _05716_ : _05715_;
  assign _05718_ = \bapg_rd.w_ptr_r [2] ? _05717_ : _05714_;
  assign _05719_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [4] : \MSYNC_1r1w.synth.nz.mem[552] [4];
  assign _05720_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [4] : \MSYNC_1r1w.synth.nz.mem[554] [4];
  assign _05721_ = \bapg_rd.w_ptr_r [1] ? _05720_ : _05719_;
  assign _05722_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [4] : \MSYNC_1r1w.synth.nz.mem[556] [4];
  assign _05723_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [4] : \MSYNC_1r1w.synth.nz.mem[558] [4];
  assign _05724_ = \bapg_rd.w_ptr_r [1] ? _05723_ : _05722_;
  assign _05725_ = \bapg_rd.w_ptr_r [2] ? _05724_ : _05721_;
  assign _05726_ = \bapg_rd.w_ptr_r [3] ? _05725_ : _05718_;
  assign _05727_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [4] : \MSYNC_1r1w.synth.nz.mem[560] [4];
  assign _05728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [4] : \MSYNC_1r1w.synth.nz.mem[562] [4];
  assign _05729_ = \bapg_rd.w_ptr_r [1] ? _05728_ : _05727_;
  assign _05730_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [4] : \MSYNC_1r1w.synth.nz.mem[564] [4];
  assign _05731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [4] : \MSYNC_1r1w.synth.nz.mem[566] [4];
  assign _05732_ = \bapg_rd.w_ptr_r [1] ? _05731_ : _05730_;
  assign _05733_ = \bapg_rd.w_ptr_r [2] ? _05732_ : _05729_;
  assign _05734_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [4] : \MSYNC_1r1w.synth.nz.mem[568] [4];
  assign _05735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [4] : \MSYNC_1r1w.synth.nz.mem[570] [4];
  assign _05736_ = \bapg_rd.w_ptr_r [1] ? _05735_ : _05734_;
  assign _05737_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [4] : \MSYNC_1r1w.synth.nz.mem[572] [4];
  assign _05738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [4] : \MSYNC_1r1w.synth.nz.mem[574] [4];
  assign _05739_ = \bapg_rd.w_ptr_r [1] ? _05738_ : _05737_;
  assign _05740_ = \bapg_rd.w_ptr_r [2] ? _05739_ : _05736_;
  assign _05741_ = \bapg_rd.w_ptr_r [3] ? _05740_ : _05733_;
  assign _05742_ = \bapg_rd.w_ptr_r [4] ? _05741_ : _05726_;
  assign _05743_ = \bapg_rd.w_ptr_r [5] ? _05742_ : _05711_;
  assign _05744_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [4] : \MSYNC_1r1w.synth.nz.mem[576] [4];
  assign _05745_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [4] : \MSYNC_1r1w.synth.nz.mem[578] [4];
  assign _05746_ = \bapg_rd.w_ptr_r [1] ? _05745_ : _05744_;
  assign _05747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [4] : \MSYNC_1r1w.synth.nz.mem[580] [4];
  assign _05748_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [4] : \MSYNC_1r1w.synth.nz.mem[582] [4];
  assign _05749_ = \bapg_rd.w_ptr_r [1] ? _05748_ : _05747_;
  assign _05750_ = \bapg_rd.w_ptr_r [2] ? _05749_ : _05746_;
  assign _05751_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [4] : \MSYNC_1r1w.synth.nz.mem[584] [4];
  assign _05752_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [4] : \MSYNC_1r1w.synth.nz.mem[586] [4];
  assign _05753_ = \bapg_rd.w_ptr_r [1] ? _05752_ : _05751_;
  assign _05754_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [4] : \MSYNC_1r1w.synth.nz.mem[588] [4];
  assign _05755_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [4] : \MSYNC_1r1w.synth.nz.mem[590] [4];
  assign _05756_ = \bapg_rd.w_ptr_r [1] ? _05755_ : _05754_;
  assign _05757_ = \bapg_rd.w_ptr_r [2] ? _05756_ : _05753_;
  assign _05758_ = \bapg_rd.w_ptr_r [3] ? _05757_ : _05750_;
  assign _05759_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [4] : \MSYNC_1r1w.synth.nz.mem[592] [4];
  assign _05760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [4] : \MSYNC_1r1w.synth.nz.mem[594] [4];
  assign _05761_ = \bapg_rd.w_ptr_r [1] ? _05760_ : _05759_;
  assign _05762_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [4] : \MSYNC_1r1w.synth.nz.mem[596] [4];
  assign _05763_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [4] : \MSYNC_1r1w.synth.nz.mem[598] [4];
  assign _05764_ = \bapg_rd.w_ptr_r [1] ? _05763_ : _05762_;
  assign _05765_ = \bapg_rd.w_ptr_r [2] ? _05764_ : _05761_;
  assign _05766_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [4] : \MSYNC_1r1w.synth.nz.mem[600] [4];
  assign _05767_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [4] : \MSYNC_1r1w.synth.nz.mem[602] [4];
  assign _05768_ = \bapg_rd.w_ptr_r [1] ? _05767_ : _05766_;
  assign _05769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [4] : \MSYNC_1r1w.synth.nz.mem[604] [4];
  assign _05770_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [4] : \MSYNC_1r1w.synth.nz.mem[606] [4];
  assign _05771_ = \bapg_rd.w_ptr_r [1] ? _05770_ : _05769_;
  assign _05772_ = \bapg_rd.w_ptr_r [2] ? _05771_ : _05768_;
  assign _05773_ = \bapg_rd.w_ptr_r [3] ? _05772_ : _05765_;
  assign _05774_ = \bapg_rd.w_ptr_r [4] ? _05773_ : _05758_;
  assign _05775_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [4] : \MSYNC_1r1w.synth.nz.mem[608] [4];
  assign _05776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [4] : \MSYNC_1r1w.synth.nz.mem[610] [4];
  assign _05777_ = \bapg_rd.w_ptr_r [1] ? _05776_ : _05775_;
  assign _05778_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [4] : \MSYNC_1r1w.synth.nz.mem[612] [4];
  assign _05779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [4] : \MSYNC_1r1w.synth.nz.mem[614] [4];
  assign _05780_ = \bapg_rd.w_ptr_r [1] ? _05779_ : _05778_;
  assign _05781_ = \bapg_rd.w_ptr_r [2] ? _05780_ : _05777_;
  assign _05782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [4] : \MSYNC_1r1w.synth.nz.mem[616] [4];
  assign _05783_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [4] : \MSYNC_1r1w.synth.nz.mem[618] [4];
  assign _05784_ = \bapg_rd.w_ptr_r [1] ? _05783_ : _05782_;
  assign _05785_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [4] : \MSYNC_1r1w.synth.nz.mem[620] [4];
  assign _05786_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [4] : \MSYNC_1r1w.synth.nz.mem[622] [4];
  assign _05787_ = \bapg_rd.w_ptr_r [1] ? _05786_ : _05785_;
  assign _05788_ = \bapg_rd.w_ptr_r [2] ? _05787_ : _05784_;
  assign _05789_ = \bapg_rd.w_ptr_r [3] ? _05788_ : _05781_;
  assign _05790_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [4] : \MSYNC_1r1w.synth.nz.mem[624] [4];
  assign _05791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [4] : \MSYNC_1r1w.synth.nz.mem[626] [4];
  assign _05792_ = \bapg_rd.w_ptr_r [1] ? _05791_ : _05790_;
  assign _05793_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [4] : \MSYNC_1r1w.synth.nz.mem[628] [4];
  assign _05794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [4] : \MSYNC_1r1w.synth.nz.mem[630] [4];
  assign _05795_ = \bapg_rd.w_ptr_r [1] ? _05794_ : _05793_;
  assign _05796_ = \bapg_rd.w_ptr_r [2] ? _05795_ : _05792_;
  assign _05797_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [4] : \MSYNC_1r1w.synth.nz.mem[632] [4];
  assign _05798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [4] : \MSYNC_1r1w.synth.nz.mem[634] [4];
  assign _05799_ = \bapg_rd.w_ptr_r [1] ? _05798_ : _05797_;
  assign _05800_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [4] : \MSYNC_1r1w.synth.nz.mem[636] [4];
  assign _05801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [4] : \MSYNC_1r1w.synth.nz.mem[638] [4];
  assign _05802_ = \bapg_rd.w_ptr_r [1] ? _05801_ : _05800_;
  assign _05803_ = \bapg_rd.w_ptr_r [2] ? _05802_ : _05799_;
  assign _05804_ = \bapg_rd.w_ptr_r [3] ? _05803_ : _05796_;
  assign _05805_ = \bapg_rd.w_ptr_r [4] ? _05804_ : _05789_;
  assign _05806_ = \bapg_rd.w_ptr_r [5] ? _05805_ : _05774_;
  assign _05807_ = \bapg_rd.w_ptr_r [6] ? _05806_ : _05743_;
  assign _05808_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [4] : \MSYNC_1r1w.synth.nz.mem[640] [4];
  assign _05809_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [4] : \MSYNC_1r1w.synth.nz.mem[642] [4];
  assign _05810_ = \bapg_rd.w_ptr_r [1] ? _05809_ : _05808_;
  assign _05811_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [4] : \MSYNC_1r1w.synth.nz.mem[644] [4];
  assign _05812_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [4] : \MSYNC_1r1w.synth.nz.mem[646] [4];
  assign _05813_ = \bapg_rd.w_ptr_r [1] ? _05812_ : _05811_;
  assign _05814_ = \bapg_rd.w_ptr_r [2] ? _05813_ : _05810_;
  assign _05815_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [4] : \MSYNC_1r1w.synth.nz.mem[648] [4];
  assign _05816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [4] : \MSYNC_1r1w.synth.nz.mem[650] [4];
  assign _05817_ = \bapg_rd.w_ptr_r [1] ? _05816_ : _05815_;
  assign _05818_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [4] : \MSYNC_1r1w.synth.nz.mem[652] [4];
  assign _05819_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [4] : \MSYNC_1r1w.synth.nz.mem[654] [4];
  assign _05820_ = \bapg_rd.w_ptr_r [1] ? _05819_ : _05818_;
  assign _05821_ = \bapg_rd.w_ptr_r [2] ? _05820_ : _05817_;
  assign _05822_ = \bapg_rd.w_ptr_r [3] ? _05821_ : _05814_;
  assign _05823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [4] : \MSYNC_1r1w.synth.nz.mem[656] [4];
  assign _05824_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [4] : \MSYNC_1r1w.synth.nz.mem[658] [4];
  assign _05825_ = \bapg_rd.w_ptr_r [1] ? _05824_ : _05823_;
  assign _05826_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [4] : \MSYNC_1r1w.synth.nz.mem[660] [4];
  assign _05827_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [4] : \MSYNC_1r1w.synth.nz.mem[662] [4];
  assign _05828_ = \bapg_rd.w_ptr_r [1] ? _05827_ : _05826_;
  assign _05829_ = \bapg_rd.w_ptr_r [2] ? _05828_ : _05825_;
  assign _05830_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [4] : \MSYNC_1r1w.synth.nz.mem[664] [4];
  assign _05831_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [4] : \MSYNC_1r1w.synth.nz.mem[666] [4];
  assign _05832_ = \bapg_rd.w_ptr_r [1] ? _05831_ : _05830_;
  assign _05833_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [4] : \MSYNC_1r1w.synth.nz.mem[668] [4];
  assign _05834_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [4] : \MSYNC_1r1w.synth.nz.mem[670] [4];
  assign _05835_ = \bapg_rd.w_ptr_r [1] ? _05834_ : _05833_;
  assign _05836_ = \bapg_rd.w_ptr_r [2] ? _05835_ : _05832_;
  assign _05837_ = \bapg_rd.w_ptr_r [3] ? _05836_ : _05829_;
  assign _05838_ = \bapg_rd.w_ptr_r [4] ? _05837_ : _05822_;
  assign _05839_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [4] : \MSYNC_1r1w.synth.nz.mem[672] [4];
  assign _05840_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [4] : \MSYNC_1r1w.synth.nz.mem[674] [4];
  assign _05841_ = \bapg_rd.w_ptr_r [1] ? _05840_ : _05839_;
  assign _05842_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [4] : \MSYNC_1r1w.synth.nz.mem[676] [4];
  assign _05843_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [4] : \MSYNC_1r1w.synth.nz.mem[678] [4];
  assign _05844_ = \bapg_rd.w_ptr_r [1] ? _05843_ : _05842_;
  assign _05845_ = \bapg_rd.w_ptr_r [2] ? _05844_ : _05841_;
  assign _05846_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [4] : \MSYNC_1r1w.synth.nz.mem[680] [4];
  assign _05847_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [4] : \MSYNC_1r1w.synth.nz.mem[682] [4];
  assign _05848_ = \bapg_rd.w_ptr_r [1] ? _05847_ : _05846_;
  assign _05849_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [4] : \MSYNC_1r1w.synth.nz.mem[684] [4];
  assign _05850_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [4] : \MSYNC_1r1w.synth.nz.mem[686] [4];
  assign _05851_ = \bapg_rd.w_ptr_r [1] ? _05850_ : _05849_;
  assign _05852_ = \bapg_rd.w_ptr_r [2] ? _05851_ : _05848_;
  assign _05853_ = \bapg_rd.w_ptr_r [3] ? _05852_ : _05845_;
  assign _05854_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [4] : \MSYNC_1r1w.synth.nz.mem[688] [4];
  assign _05855_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [4] : \MSYNC_1r1w.synth.nz.mem[690] [4];
  assign _05856_ = \bapg_rd.w_ptr_r [1] ? _05855_ : _05854_;
  assign _05857_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [4] : \MSYNC_1r1w.synth.nz.mem[692] [4];
  assign _05858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [4] : \MSYNC_1r1w.synth.nz.mem[694] [4];
  assign _05859_ = \bapg_rd.w_ptr_r [1] ? _05858_ : _05857_;
  assign _05860_ = \bapg_rd.w_ptr_r [2] ? _05859_ : _05856_;
  assign _05861_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [4] : \MSYNC_1r1w.synth.nz.mem[696] [4];
  assign _05862_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [4] : \MSYNC_1r1w.synth.nz.mem[698] [4];
  assign _05863_ = \bapg_rd.w_ptr_r [1] ? _05862_ : _05861_;
  assign _05864_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [4] : \MSYNC_1r1w.synth.nz.mem[700] [4];
  assign _05865_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [4] : \MSYNC_1r1w.synth.nz.mem[702] [4];
  assign _05866_ = \bapg_rd.w_ptr_r [1] ? _05865_ : _05864_;
  assign _05867_ = \bapg_rd.w_ptr_r [2] ? _05866_ : _05863_;
  assign _05868_ = \bapg_rd.w_ptr_r [3] ? _05867_ : _05860_;
  assign _05869_ = \bapg_rd.w_ptr_r [4] ? _05868_ : _05853_;
  assign _05870_ = \bapg_rd.w_ptr_r [5] ? _05869_ : _05838_;
  assign _05871_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [4] : \MSYNC_1r1w.synth.nz.mem[704] [4];
  assign _05872_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [4] : \MSYNC_1r1w.synth.nz.mem[706] [4];
  assign _05873_ = \bapg_rd.w_ptr_r [1] ? _05872_ : _05871_;
  assign _05874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [4] : \MSYNC_1r1w.synth.nz.mem[708] [4];
  assign _05875_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [4] : \MSYNC_1r1w.synth.nz.mem[710] [4];
  assign _05876_ = \bapg_rd.w_ptr_r [1] ? _05875_ : _05874_;
  assign _05877_ = \bapg_rd.w_ptr_r [2] ? _05876_ : _05873_;
  assign _05878_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [4] : \MSYNC_1r1w.synth.nz.mem[712] [4];
  assign _05879_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [4] : \MSYNC_1r1w.synth.nz.mem[714] [4];
  assign _05880_ = \bapg_rd.w_ptr_r [1] ? _05879_ : _05878_;
  assign _05881_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [4] : \MSYNC_1r1w.synth.nz.mem[716] [4];
  assign _05882_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [4] : \MSYNC_1r1w.synth.nz.mem[718] [4];
  assign _05883_ = \bapg_rd.w_ptr_r [1] ? _05882_ : _05881_;
  assign _05884_ = \bapg_rd.w_ptr_r [2] ? _05883_ : _05880_;
  assign _05885_ = \bapg_rd.w_ptr_r [3] ? _05884_ : _05877_;
  assign _05886_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [4] : \MSYNC_1r1w.synth.nz.mem[720] [4];
  assign _05887_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [4] : \MSYNC_1r1w.synth.nz.mem[722] [4];
  assign _05888_ = \bapg_rd.w_ptr_r [1] ? _05887_ : _05886_;
  assign _05889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [4] : \MSYNC_1r1w.synth.nz.mem[724] [4];
  assign _05890_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [4] : \MSYNC_1r1w.synth.nz.mem[726] [4];
  assign _05891_ = \bapg_rd.w_ptr_r [1] ? _05890_ : _05889_;
  assign _05892_ = \bapg_rd.w_ptr_r [2] ? _05891_ : _05888_;
  assign _05893_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [4] : \MSYNC_1r1w.synth.nz.mem[728] [4];
  assign _05894_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [4] : \MSYNC_1r1w.synth.nz.mem[730] [4];
  assign _05895_ = \bapg_rd.w_ptr_r [1] ? _05894_ : _05893_;
  assign _05896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [4] : \MSYNC_1r1w.synth.nz.mem[732] [4];
  assign _05897_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [4] : \MSYNC_1r1w.synth.nz.mem[734] [4];
  assign _05898_ = \bapg_rd.w_ptr_r [1] ? _05897_ : _05896_;
  assign _05899_ = \bapg_rd.w_ptr_r [2] ? _05898_ : _05895_;
  assign _05900_ = \bapg_rd.w_ptr_r [3] ? _05899_ : _05892_;
  assign _05901_ = \bapg_rd.w_ptr_r [4] ? _05900_ : _05885_;
  assign _05902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [4] : \MSYNC_1r1w.synth.nz.mem[736] [4];
  assign _05903_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [4] : \MSYNC_1r1w.synth.nz.mem[738] [4];
  assign _05904_ = \bapg_rd.w_ptr_r [1] ? _05903_ : _05902_;
  assign _05905_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [4] : \MSYNC_1r1w.synth.nz.mem[740] [4];
  assign _05906_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [4] : \MSYNC_1r1w.synth.nz.mem[742] [4];
  assign _05907_ = \bapg_rd.w_ptr_r [1] ? _05906_ : _05905_;
  assign _05908_ = \bapg_rd.w_ptr_r [2] ? _05907_ : _05904_;
  assign _05909_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [4] : \MSYNC_1r1w.synth.nz.mem[744] [4];
  assign _05910_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [4] : \MSYNC_1r1w.synth.nz.mem[746] [4];
  assign _05911_ = \bapg_rd.w_ptr_r [1] ? _05910_ : _05909_;
  assign _05912_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [4] : \MSYNC_1r1w.synth.nz.mem[748] [4];
  assign _05913_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [4] : \MSYNC_1r1w.synth.nz.mem[750] [4];
  assign _05914_ = \bapg_rd.w_ptr_r [1] ? _05913_ : _05912_;
  assign _05915_ = \bapg_rd.w_ptr_r [2] ? _05914_ : _05911_;
  assign _05916_ = \bapg_rd.w_ptr_r [3] ? _05915_ : _05908_;
  assign _05917_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [4] : \MSYNC_1r1w.synth.nz.mem[752] [4];
  assign _05918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [4] : \MSYNC_1r1w.synth.nz.mem[754] [4];
  assign _05919_ = \bapg_rd.w_ptr_r [1] ? _05918_ : _05917_;
  assign _05920_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [4] : \MSYNC_1r1w.synth.nz.mem[756] [4];
  assign _05921_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [4] : \MSYNC_1r1w.synth.nz.mem[758] [4];
  assign _05922_ = \bapg_rd.w_ptr_r [1] ? _05921_ : _05920_;
  assign _05923_ = \bapg_rd.w_ptr_r [2] ? _05922_ : _05919_;
  assign _05924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [4] : \MSYNC_1r1w.synth.nz.mem[760] [4];
  assign _05925_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [4] : \MSYNC_1r1w.synth.nz.mem[762] [4];
  assign _05926_ = \bapg_rd.w_ptr_r [1] ? _05925_ : _05924_;
  assign _05927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [4] : \MSYNC_1r1w.synth.nz.mem[764] [4];
  assign _05928_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [4] : \MSYNC_1r1w.synth.nz.mem[766] [4];
  assign _05929_ = \bapg_rd.w_ptr_r [1] ? _05928_ : _05927_;
  assign _05930_ = \bapg_rd.w_ptr_r [2] ? _05929_ : _05926_;
  assign _05931_ = \bapg_rd.w_ptr_r [3] ? _05930_ : _05923_;
  assign _05932_ = \bapg_rd.w_ptr_r [4] ? _05931_ : _05916_;
  assign _05933_ = \bapg_rd.w_ptr_r [5] ? _05932_ : _05901_;
  assign _05934_ = \bapg_rd.w_ptr_r [6] ? _05933_ : _05870_;
  assign _05935_ = \bapg_rd.w_ptr_r [7] ? _05934_ : _05807_;
  assign _05936_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [4] : \MSYNC_1r1w.synth.nz.mem[768] [4];
  assign _05937_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [4] : \MSYNC_1r1w.synth.nz.mem[770] [4];
  assign _05938_ = \bapg_rd.w_ptr_r [1] ? _05937_ : _05936_;
  assign _05939_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [4] : \MSYNC_1r1w.synth.nz.mem[772] [4];
  assign _05940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [4] : \MSYNC_1r1w.synth.nz.mem[774] [4];
  assign _05941_ = \bapg_rd.w_ptr_r [1] ? _05940_ : _05939_;
  assign _05942_ = \bapg_rd.w_ptr_r [2] ? _05941_ : _05938_;
  assign _05943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [4] : \MSYNC_1r1w.synth.nz.mem[776] [4];
  assign _05944_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [4] : \MSYNC_1r1w.synth.nz.mem[778] [4];
  assign _05945_ = \bapg_rd.w_ptr_r [1] ? _05944_ : _05943_;
  assign _05946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [4] : \MSYNC_1r1w.synth.nz.mem[780] [4];
  assign _05947_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [4] : \MSYNC_1r1w.synth.nz.mem[782] [4];
  assign _05948_ = \bapg_rd.w_ptr_r [1] ? _05947_ : _05946_;
  assign _05949_ = \bapg_rd.w_ptr_r [2] ? _05948_ : _05945_;
  assign _05950_ = \bapg_rd.w_ptr_r [3] ? _05949_ : _05942_;
  assign _05951_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [4] : \MSYNC_1r1w.synth.nz.mem[784] [4];
  assign _05952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [4] : \MSYNC_1r1w.synth.nz.mem[786] [4];
  assign _05953_ = \bapg_rd.w_ptr_r [1] ? _05952_ : _05951_;
  assign _05954_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [4] : \MSYNC_1r1w.synth.nz.mem[788] [4];
  assign _05955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [4] : \MSYNC_1r1w.synth.nz.mem[790] [4];
  assign _05956_ = \bapg_rd.w_ptr_r [1] ? _05955_ : _05954_;
  assign _05957_ = \bapg_rd.w_ptr_r [2] ? _05956_ : _05953_;
  assign _05958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [4] : \MSYNC_1r1w.synth.nz.mem[792] [4];
  assign _05959_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [4] : \MSYNC_1r1w.synth.nz.mem[794] [4];
  assign _05960_ = \bapg_rd.w_ptr_r [1] ? _05959_ : _05958_;
  assign _05961_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [4] : \MSYNC_1r1w.synth.nz.mem[796] [4];
  assign _05962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [4] : \MSYNC_1r1w.synth.nz.mem[798] [4];
  assign _05963_ = \bapg_rd.w_ptr_r [1] ? _05962_ : _05961_;
  assign _05964_ = \bapg_rd.w_ptr_r [2] ? _05963_ : _05960_;
  assign _05965_ = \bapg_rd.w_ptr_r [3] ? _05964_ : _05957_;
  assign _05966_ = \bapg_rd.w_ptr_r [4] ? _05965_ : _05950_;
  assign _05967_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [4] : \MSYNC_1r1w.synth.nz.mem[800] [4];
  assign _05968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [4] : \MSYNC_1r1w.synth.nz.mem[802] [4];
  assign _05969_ = \bapg_rd.w_ptr_r [1] ? _05968_ : _05967_;
  assign _05970_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [4] : \MSYNC_1r1w.synth.nz.mem[804] [4];
  assign _05971_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [4] : \MSYNC_1r1w.synth.nz.mem[806] [4];
  assign _05972_ = \bapg_rd.w_ptr_r [1] ? _05971_ : _05970_;
  assign _05973_ = \bapg_rd.w_ptr_r [2] ? _05972_ : _05969_;
  assign _05974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [4] : \MSYNC_1r1w.synth.nz.mem[808] [4];
  assign _05975_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [4] : \MSYNC_1r1w.synth.nz.mem[810] [4];
  assign _05976_ = \bapg_rd.w_ptr_r [1] ? _05975_ : _05974_;
  assign _05977_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [4] : \MSYNC_1r1w.synth.nz.mem[812] [4];
  assign _05978_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [4] : \MSYNC_1r1w.synth.nz.mem[814] [4];
  assign _05979_ = \bapg_rd.w_ptr_r [1] ? _05978_ : _05977_;
  assign _05980_ = \bapg_rd.w_ptr_r [2] ? _05979_ : _05976_;
  assign _05981_ = \bapg_rd.w_ptr_r [3] ? _05980_ : _05973_;
  assign _05982_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [4] : \MSYNC_1r1w.synth.nz.mem[816] [4];
  assign _05983_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [4] : \MSYNC_1r1w.synth.nz.mem[818] [4];
  assign _05984_ = \bapg_rd.w_ptr_r [1] ? _05983_ : _05982_;
  assign _05985_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [4] : \MSYNC_1r1w.synth.nz.mem[820] [4];
  assign _05986_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [4] : \MSYNC_1r1w.synth.nz.mem[822] [4];
  assign _05987_ = \bapg_rd.w_ptr_r [1] ? _05986_ : _05985_;
  assign _05988_ = \bapg_rd.w_ptr_r [2] ? _05987_ : _05984_;
  assign _05989_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [4] : \MSYNC_1r1w.synth.nz.mem[824] [4];
  assign _05990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [4] : \MSYNC_1r1w.synth.nz.mem[826] [4];
  assign _05991_ = \bapg_rd.w_ptr_r [1] ? _05990_ : _05989_;
  assign _05992_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [4] : \MSYNC_1r1w.synth.nz.mem[828] [4];
  assign _05993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [4] : \MSYNC_1r1w.synth.nz.mem[830] [4];
  assign _05994_ = \bapg_rd.w_ptr_r [1] ? _05993_ : _05992_;
  assign _05995_ = \bapg_rd.w_ptr_r [2] ? _05994_ : _05991_;
  assign _05996_ = \bapg_rd.w_ptr_r [3] ? _05995_ : _05988_;
  assign _05997_ = \bapg_rd.w_ptr_r [4] ? _05996_ : _05981_;
  assign _05998_ = \bapg_rd.w_ptr_r [5] ? _05997_ : _05966_;
  assign _05999_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [4] : \MSYNC_1r1w.synth.nz.mem[832] [4];
  assign _06000_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [4] : \MSYNC_1r1w.synth.nz.mem[834] [4];
  assign _06001_ = \bapg_rd.w_ptr_r [1] ? _06000_ : _05999_;
  assign _06002_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [4] : \MSYNC_1r1w.synth.nz.mem[836] [4];
  assign _06003_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [4] : \MSYNC_1r1w.synth.nz.mem[838] [4];
  assign _06004_ = \bapg_rd.w_ptr_r [1] ? _06003_ : _06002_;
  assign _06005_ = \bapg_rd.w_ptr_r [2] ? _06004_ : _06001_;
  assign _06006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [4] : \MSYNC_1r1w.synth.nz.mem[840] [4];
  assign _06007_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [4] : \MSYNC_1r1w.synth.nz.mem[842] [4];
  assign _06008_ = \bapg_rd.w_ptr_r [1] ? _06007_ : _06006_;
  assign _06009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [4] : \MSYNC_1r1w.synth.nz.mem[844] [4];
  assign _06010_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [4] : \MSYNC_1r1w.synth.nz.mem[846] [4];
  assign _06011_ = \bapg_rd.w_ptr_r [1] ? _06010_ : _06009_;
  assign _06012_ = \bapg_rd.w_ptr_r [2] ? _06011_ : _06008_;
  assign _06013_ = \bapg_rd.w_ptr_r [3] ? _06012_ : _06005_;
  assign _06014_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [4] : \MSYNC_1r1w.synth.nz.mem[848] [4];
  assign _06015_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [4] : \MSYNC_1r1w.synth.nz.mem[850] [4];
  assign _06016_ = \bapg_rd.w_ptr_r [1] ? _06015_ : _06014_;
  assign _06017_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [4] : \MSYNC_1r1w.synth.nz.mem[852] [4];
  assign _06018_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [4] : \MSYNC_1r1w.synth.nz.mem[854] [4];
  assign _06019_ = \bapg_rd.w_ptr_r [1] ? _06018_ : _06017_;
  assign _06020_ = \bapg_rd.w_ptr_r [2] ? _06019_ : _06016_;
  assign _06021_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [4] : \MSYNC_1r1w.synth.nz.mem[856] [4];
  assign _06022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [4] : \MSYNC_1r1w.synth.nz.mem[858] [4];
  assign _06023_ = \bapg_rd.w_ptr_r [1] ? _06022_ : _06021_;
  assign _06024_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [4] : \MSYNC_1r1w.synth.nz.mem[860] [4];
  assign _06025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [4] : \MSYNC_1r1w.synth.nz.mem[862] [4];
  assign _06026_ = \bapg_rd.w_ptr_r [1] ? _06025_ : _06024_;
  assign _06027_ = \bapg_rd.w_ptr_r [2] ? _06026_ : _06023_;
  assign _06028_ = \bapg_rd.w_ptr_r [3] ? _06027_ : _06020_;
  assign _06029_ = \bapg_rd.w_ptr_r [4] ? _06028_ : _06013_;
  assign _06030_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [4] : \MSYNC_1r1w.synth.nz.mem[864] [4];
  assign _06031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [4] : \MSYNC_1r1w.synth.nz.mem[866] [4];
  assign _06032_ = \bapg_rd.w_ptr_r [1] ? _06031_ : _06030_;
  assign _06033_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [4] : \MSYNC_1r1w.synth.nz.mem[868] [4];
  assign _06034_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [4] : \MSYNC_1r1w.synth.nz.mem[870] [4];
  assign _06035_ = \bapg_rd.w_ptr_r [1] ? _06034_ : _06033_;
  assign _06036_ = \bapg_rd.w_ptr_r [2] ? _06035_ : _06032_;
  assign _06037_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [4] : \MSYNC_1r1w.synth.nz.mem[872] [4];
  assign _06038_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [4] : \MSYNC_1r1w.synth.nz.mem[874] [4];
  assign _06039_ = \bapg_rd.w_ptr_r [1] ? _06038_ : _06037_;
  assign _06040_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [4] : \MSYNC_1r1w.synth.nz.mem[876] [4];
  assign _06041_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [4] : \MSYNC_1r1w.synth.nz.mem[878] [4];
  assign _06042_ = \bapg_rd.w_ptr_r [1] ? _06041_ : _06040_;
  assign _06043_ = \bapg_rd.w_ptr_r [2] ? _06042_ : _06039_;
  assign _06044_ = \bapg_rd.w_ptr_r [3] ? _06043_ : _06036_;
  assign _06045_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [4] : \MSYNC_1r1w.synth.nz.mem[880] [4];
  assign _06046_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [4] : \MSYNC_1r1w.synth.nz.mem[882] [4];
  assign _06047_ = \bapg_rd.w_ptr_r [1] ? _06046_ : _06045_;
  assign _06048_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [4] : \MSYNC_1r1w.synth.nz.mem[884] [4];
  assign _06049_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [4] : \MSYNC_1r1w.synth.nz.mem[886] [4];
  assign _06050_ = \bapg_rd.w_ptr_r [1] ? _06049_ : _06048_;
  assign _06051_ = \bapg_rd.w_ptr_r [2] ? _06050_ : _06047_;
  assign _06052_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [4] : \MSYNC_1r1w.synth.nz.mem[888] [4];
  assign _06053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [4] : \MSYNC_1r1w.synth.nz.mem[890] [4];
  assign _06054_ = \bapg_rd.w_ptr_r [1] ? _06053_ : _06052_;
  assign _06055_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [4] : \MSYNC_1r1w.synth.nz.mem[892] [4];
  assign _06056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [4] : \MSYNC_1r1w.synth.nz.mem[894] [4];
  assign _06057_ = \bapg_rd.w_ptr_r [1] ? _06056_ : _06055_;
  assign _06058_ = \bapg_rd.w_ptr_r [2] ? _06057_ : _06054_;
  assign _06059_ = \bapg_rd.w_ptr_r [3] ? _06058_ : _06051_;
  assign _06060_ = \bapg_rd.w_ptr_r [4] ? _06059_ : _06044_;
  assign _06061_ = \bapg_rd.w_ptr_r [5] ? _06060_ : _06029_;
  assign _06062_ = \bapg_rd.w_ptr_r [6] ? _06061_ : _05998_;
  assign _06063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [4] : \MSYNC_1r1w.synth.nz.mem[896] [4];
  assign _06064_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [4] : \MSYNC_1r1w.synth.nz.mem[898] [4];
  assign _06065_ = \bapg_rd.w_ptr_r [1] ? _06064_ : _06063_;
  assign _06066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [4] : \MSYNC_1r1w.synth.nz.mem[900] [4];
  assign _06067_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [4] : \MSYNC_1r1w.synth.nz.mem[902] [4];
  assign _06068_ = \bapg_rd.w_ptr_r [1] ? _06067_ : _06066_;
  assign _06069_ = \bapg_rd.w_ptr_r [2] ? _06068_ : _06065_;
  assign _06070_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [4] : \MSYNC_1r1w.synth.nz.mem[904] [4];
  assign _06071_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [4] : \MSYNC_1r1w.synth.nz.mem[906] [4];
  assign _06072_ = \bapg_rd.w_ptr_r [1] ? _06071_ : _06070_;
  assign _06073_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [4] : \MSYNC_1r1w.synth.nz.mem[908] [4];
  assign _06074_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [4] : \MSYNC_1r1w.synth.nz.mem[910] [4];
  assign _06075_ = \bapg_rd.w_ptr_r [1] ? _06074_ : _06073_;
  assign _06076_ = \bapg_rd.w_ptr_r [2] ? _06075_ : _06072_;
  assign _06077_ = \bapg_rd.w_ptr_r [3] ? _06076_ : _06069_;
  assign _06078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [4] : \MSYNC_1r1w.synth.nz.mem[912] [4];
  assign _06079_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [4] : \MSYNC_1r1w.synth.nz.mem[914] [4];
  assign _06080_ = \bapg_rd.w_ptr_r [1] ? _06079_ : _06078_;
  assign _06081_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [4] : \MSYNC_1r1w.synth.nz.mem[916] [4];
  assign _06082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [4] : \MSYNC_1r1w.synth.nz.mem[918] [4];
  assign _06083_ = \bapg_rd.w_ptr_r [1] ? _06082_ : _06081_;
  assign _06084_ = \bapg_rd.w_ptr_r [2] ? _06083_ : _06080_;
  assign _06085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [4] : \MSYNC_1r1w.synth.nz.mem[920] [4];
  assign _06086_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [4] : \MSYNC_1r1w.synth.nz.mem[922] [4];
  assign _06087_ = \bapg_rd.w_ptr_r [1] ? _06086_ : _06085_;
  assign _06088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [4] : \MSYNC_1r1w.synth.nz.mem[924] [4];
  assign _06089_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [4] : \MSYNC_1r1w.synth.nz.mem[926] [4];
  assign _06090_ = \bapg_rd.w_ptr_r [1] ? _06089_ : _06088_;
  assign _06091_ = \bapg_rd.w_ptr_r [2] ? _06090_ : _06087_;
  assign _06092_ = \bapg_rd.w_ptr_r [3] ? _06091_ : _06084_;
  assign _06093_ = \bapg_rd.w_ptr_r [4] ? _06092_ : _06077_;
  assign _06094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [4] : \MSYNC_1r1w.synth.nz.mem[928] [4];
  assign _06095_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [4] : \MSYNC_1r1w.synth.nz.mem[930] [4];
  assign _06096_ = \bapg_rd.w_ptr_r [1] ? _06095_ : _06094_;
  assign _06097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [4] : \MSYNC_1r1w.synth.nz.mem[932] [4];
  assign _06098_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [4] : \MSYNC_1r1w.synth.nz.mem[934] [4];
  assign _06099_ = \bapg_rd.w_ptr_r [1] ? _06098_ : _06097_;
  assign _06100_ = \bapg_rd.w_ptr_r [2] ? _06099_ : _06096_;
  assign _06101_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [4] : \MSYNC_1r1w.synth.nz.mem[936] [4];
  assign _06102_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [4] : \MSYNC_1r1w.synth.nz.mem[938] [4];
  assign _06103_ = \bapg_rd.w_ptr_r [1] ? _06102_ : _06101_;
  assign _06104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [4] : \MSYNC_1r1w.synth.nz.mem[940] [4];
  assign _06105_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [4] : \MSYNC_1r1w.synth.nz.mem[942] [4];
  assign _06106_ = \bapg_rd.w_ptr_r [1] ? _06105_ : _06104_;
  assign _06107_ = \bapg_rd.w_ptr_r [2] ? _06106_ : _06103_;
  assign _06108_ = \bapg_rd.w_ptr_r [3] ? _06107_ : _06100_;
  assign _06109_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [4] : \MSYNC_1r1w.synth.nz.mem[944] [4];
  assign _06110_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [4] : \MSYNC_1r1w.synth.nz.mem[946] [4];
  assign _06111_ = \bapg_rd.w_ptr_r [1] ? _06110_ : _06109_;
  assign _06112_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [4] : \MSYNC_1r1w.synth.nz.mem[948] [4];
  assign _06113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [4] : \MSYNC_1r1w.synth.nz.mem[950] [4];
  assign _06114_ = \bapg_rd.w_ptr_r [1] ? _06113_ : _06112_;
  assign _06115_ = \bapg_rd.w_ptr_r [2] ? _06114_ : _06111_;
  assign _06116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [4] : \MSYNC_1r1w.synth.nz.mem[952] [4];
  assign _06117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [4] : \MSYNC_1r1w.synth.nz.mem[954] [4];
  assign _06118_ = \bapg_rd.w_ptr_r [1] ? _06117_ : _06116_;
  assign _06119_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [4] : \MSYNC_1r1w.synth.nz.mem[956] [4];
  assign _06120_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [4] : \MSYNC_1r1w.synth.nz.mem[958] [4];
  assign _06121_ = \bapg_rd.w_ptr_r [1] ? _06120_ : _06119_;
  assign _06122_ = \bapg_rd.w_ptr_r [2] ? _06121_ : _06118_;
  assign _06123_ = \bapg_rd.w_ptr_r [3] ? _06122_ : _06115_;
  assign _06124_ = \bapg_rd.w_ptr_r [4] ? _06123_ : _06108_;
  assign _06125_ = \bapg_rd.w_ptr_r [5] ? _06124_ : _06093_;
  assign _06126_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [4] : \MSYNC_1r1w.synth.nz.mem[960] [4];
  assign _06127_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [4] : \MSYNC_1r1w.synth.nz.mem[962] [4];
  assign _06128_ = \bapg_rd.w_ptr_r [1] ? _06127_ : _06126_;
  assign _06129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [4] : \MSYNC_1r1w.synth.nz.mem[964] [4];
  assign _06130_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [4] : \MSYNC_1r1w.synth.nz.mem[966] [4];
  assign _06131_ = \bapg_rd.w_ptr_r [1] ? _06130_ : _06129_;
  assign _06132_ = \bapg_rd.w_ptr_r [2] ? _06131_ : _06128_;
  assign _06133_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [4] : \MSYNC_1r1w.synth.nz.mem[968] [4];
  assign _06134_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [4] : \MSYNC_1r1w.synth.nz.mem[970] [4];
  assign _06135_ = \bapg_rd.w_ptr_r [1] ? _06134_ : _06133_;
  assign _06136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [4] : \MSYNC_1r1w.synth.nz.mem[972] [4];
  assign _06137_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [4] : \MSYNC_1r1w.synth.nz.mem[974] [4];
  assign _06138_ = \bapg_rd.w_ptr_r [1] ? _06137_ : _06136_;
  assign _06139_ = \bapg_rd.w_ptr_r [2] ? _06138_ : _06135_;
  assign _06140_ = \bapg_rd.w_ptr_r [3] ? _06139_ : _06132_;
  assign _06141_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [4] : \MSYNC_1r1w.synth.nz.mem[976] [4];
  assign _06142_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [4] : \MSYNC_1r1w.synth.nz.mem[978] [4];
  assign _06143_ = \bapg_rd.w_ptr_r [1] ? _06142_ : _06141_;
  assign _06144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [4] : \MSYNC_1r1w.synth.nz.mem[980] [4];
  assign _06145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [4] : \MSYNC_1r1w.synth.nz.mem[982] [4];
  assign _06146_ = \bapg_rd.w_ptr_r [1] ? _06145_ : _06144_;
  assign _06147_ = \bapg_rd.w_ptr_r [2] ? _06146_ : _06143_;
  assign _06148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [4] : \MSYNC_1r1w.synth.nz.mem[984] [4];
  assign _06149_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [4] : \MSYNC_1r1w.synth.nz.mem[986] [4];
  assign _06150_ = \bapg_rd.w_ptr_r [1] ? _06149_ : _06148_;
  assign _06151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [4] : \MSYNC_1r1w.synth.nz.mem[988] [4];
  assign _06152_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [4] : \MSYNC_1r1w.synth.nz.mem[990] [4];
  assign _06153_ = \bapg_rd.w_ptr_r [1] ? _06152_ : _06151_;
  assign _06154_ = \bapg_rd.w_ptr_r [2] ? _06153_ : _06150_;
  assign _06155_ = \bapg_rd.w_ptr_r [3] ? _06154_ : _06147_;
  assign _06156_ = \bapg_rd.w_ptr_r [4] ? _06155_ : _06140_;
  assign _06157_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [4] : \MSYNC_1r1w.synth.nz.mem[992] [4];
  assign _06158_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [4] : \MSYNC_1r1w.synth.nz.mem[994] [4];
  assign _06159_ = \bapg_rd.w_ptr_r [1] ? _06158_ : _06157_;
  assign _06160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [4] : \MSYNC_1r1w.synth.nz.mem[996] [4];
  assign _06161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [4] : \MSYNC_1r1w.synth.nz.mem[998] [4];
  assign _06162_ = \bapg_rd.w_ptr_r [1] ? _06161_ : _06160_;
  assign _06163_ = \bapg_rd.w_ptr_r [2] ? _06162_ : _06159_;
  assign _06164_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [4] : \MSYNC_1r1w.synth.nz.mem[1000] [4];
  assign _06165_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [4] : \MSYNC_1r1w.synth.nz.mem[1002] [4];
  assign _06166_ = \bapg_rd.w_ptr_r [1] ? _06165_ : _06164_;
  assign _06167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [4] : \MSYNC_1r1w.synth.nz.mem[1004] [4];
  assign _06168_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [4] : \MSYNC_1r1w.synth.nz.mem[1006] [4];
  assign _06169_ = \bapg_rd.w_ptr_r [1] ? _06168_ : _06167_;
  assign _06170_ = \bapg_rd.w_ptr_r [2] ? _06169_ : _06166_;
  assign _06171_ = \bapg_rd.w_ptr_r [3] ? _06170_ : _06163_;
  assign _06172_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [4] : \MSYNC_1r1w.synth.nz.mem[1008] [4];
  assign _06173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [4] : \MSYNC_1r1w.synth.nz.mem[1010] [4];
  assign _06174_ = \bapg_rd.w_ptr_r [1] ? _06173_ : _06172_;
  assign _06175_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [4] : \MSYNC_1r1w.synth.nz.mem[1012] [4];
  assign _06176_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [4] : \MSYNC_1r1w.synth.nz.mem[1014] [4];
  assign _06177_ = \bapg_rd.w_ptr_r [1] ? _06176_ : _06175_;
  assign _06178_ = \bapg_rd.w_ptr_r [2] ? _06177_ : _06174_;
  assign _06179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [4] : \MSYNC_1r1w.synth.nz.mem[1016] [4];
  assign _06180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [4] : \MSYNC_1r1w.synth.nz.mem[1018] [4];
  assign _06181_ = \bapg_rd.w_ptr_r [1] ? _06180_ : _06179_;
  assign _06182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [4] : \MSYNC_1r1w.synth.nz.mem[1020] [4];
  assign _06183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [4] : \MSYNC_1r1w.synth.nz.mem[1022] [4];
  assign _06184_ = \bapg_rd.w_ptr_r [1] ? _06183_ : _06182_;
  assign _06185_ = \bapg_rd.w_ptr_r [2] ? _06184_ : _06181_;
  assign _06186_ = \bapg_rd.w_ptr_r [3] ? _06185_ : _06178_;
  assign _06187_ = \bapg_rd.w_ptr_r [4] ? _06186_ : _06171_;
  assign _06188_ = \bapg_rd.w_ptr_r [5] ? _06187_ : _06156_;
  assign _06189_ = \bapg_rd.w_ptr_r [6] ? _06188_ : _06125_;
  assign _06190_ = \bapg_rd.w_ptr_r [7] ? _06189_ : _06062_;
  assign _06191_ = \bapg_rd.w_ptr_r [8] ? _06190_ : _05935_;
  assign r_data_o[4] = \bapg_rd.w_ptr_r [9] ? _06191_ : _05680_;
  assign _06192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [5] : \MSYNC_1r1w.synth.nz.mem[0] [5];
  assign _06193_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [5] : \MSYNC_1r1w.synth.nz.mem[2] [5];
  assign _06194_ = \bapg_rd.w_ptr_r [1] ? _06193_ : _06192_;
  assign _06195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [5] : \MSYNC_1r1w.synth.nz.mem[4] [5];
  assign _06196_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [5] : \MSYNC_1r1w.synth.nz.mem[6] [5];
  assign _06197_ = \bapg_rd.w_ptr_r [1] ? _06196_ : _06195_;
  assign _06198_ = \bapg_rd.w_ptr_r [2] ? _06197_ : _06194_;
  assign _06199_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [5] : \MSYNC_1r1w.synth.nz.mem[8] [5];
  assign _06200_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [5] : \MSYNC_1r1w.synth.nz.mem[10] [5];
  assign _06201_ = \bapg_rd.w_ptr_r [1] ? _06200_ : _06199_;
  assign _06202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [5] : \MSYNC_1r1w.synth.nz.mem[12] [5];
  assign _06203_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [5] : \MSYNC_1r1w.synth.nz.mem[14] [5];
  assign _06204_ = \bapg_rd.w_ptr_r [1] ? _06203_ : _06202_;
  assign _06205_ = \bapg_rd.w_ptr_r [2] ? _06204_ : _06201_;
  assign _06206_ = \bapg_rd.w_ptr_r [3] ? _06205_ : _06198_;
  assign _06207_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [5] : \MSYNC_1r1w.synth.nz.mem[16] [5];
  assign _06208_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [5] : \MSYNC_1r1w.synth.nz.mem[18] [5];
  assign _06209_ = \bapg_rd.w_ptr_r [1] ? _06208_ : _06207_;
  assign _06210_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [5] : \MSYNC_1r1w.synth.nz.mem[20] [5];
  assign _06211_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [5] : \MSYNC_1r1w.synth.nz.mem[22] [5];
  assign _06212_ = \bapg_rd.w_ptr_r [1] ? _06211_ : _06210_;
  assign _06213_ = \bapg_rd.w_ptr_r [2] ? _06212_ : _06209_;
  assign _06214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [5] : \MSYNC_1r1w.synth.nz.mem[24] [5];
  assign _06215_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [5] : \MSYNC_1r1w.synth.nz.mem[26] [5];
  assign _06216_ = \bapg_rd.w_ptr_r [1] ? _06215_ : _06214_;
  assign _06217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [5] : \MSYNC_1r1w.synth.nz.mem[28] [5];
  assign _06218_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [5] : \MSYNC_1r1w.synth.nz.mem[30] [5];
  assign _06219_ = \bapg_rd.w_ptr_r [1] ? _06218_ : _06217_;
  assign _06220_ = \bapg_rd.w_ptr_r [2] ? _06219_ : _06216_;
  assign _06221_ = \bapg_rd.w_ptr_r [3] ? _06220_ : _06213_;
  assign _06222_ = \bapg_rd.w_ptr_r [4] ? _06221_ : _06206_;
  assign _06223_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [5] : \MSYNC_1r1w.synth.nz.mem[32] [5];
  assign _06224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [5] : \MSYNC_1r1w.synth.nz.mem[34] [5];
  assign _06225_ = \bapg_rd.w_ptr_r [1] ? _06224_ : _06223_;
  assign _06226_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [5] : \MSYNC_1r1w.synth.nz.mem[36] [5];
  assign _06227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [5] : \MSYNC_1r1w.synth.nz.mem[38] [5];
  assign _06228_ = \bapg_rd.w_ptr_r [1] ? _06227_ : _06226_;
  assign _06229_ = \bapg_rd.w_ptr_r [2] ? _06228_ : _06225_;
  assign _06230_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [5] : \MSYNC_1r1w.synth.nz.mem[40] [5];
  assign _06231_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [5] : \MSYNC_1r1w.synth.nz.mem[42] [5];
  assign _06232_ = \bapg_rd.w_ptr_r [1] ? _06231_ : _06230_;
  assign _06233_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [5] : \MSYNC_1r1w.synth.nz.mem[44] [5];
  assign _06234_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [5] : \MSYNC_1r1w.synth.nz.mem[46] [5];
  assign _06235_ = \bapg_rd.w_ptr_r [1] ? _06234_ : _06233_;
  assign _06236_ = \bapg_rd.w_ptr_r [2] ? _06235_ : _06232_;
  assign _06237_ = \bapg_rd.w_ptr_r [3] ? _06236_ : _06229_;
  assign _06238_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [5] : \MSYNC_1r1w.synth.nz.mem[48] [5];
  assign _06239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [5] : \MSYNC_1r1w.synth.nz.mem[50] [5];
  assign _06240_ = \bapg_rd.w_ptr_r [1] ? _06239_ : _06238_;
  assign _06241_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [5] : \MSYNC_1r1w.synth.nz.mem[52] [5];
  assign _06242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [5] : \MSYNC_1r1w.synth.nz.mem[54] [5];
  assign _06243_ = \bapg_rd.w_ptr_r [1] ? _06242_ : _06241_;
  assign _06244_ = \bapg_rd.w_ptr_r [2] ? _06243_ : _06240_;
  assign _06245_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [5] : \MSYNC_1r1w.synth.nz.mem[56] [5];
  assign _06246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [5] : \MSYNC_1r1w.synth.nz.mem[58] [5];
  assign _06247_ = \bapg_rd.w_ptr_r [1] ? _06246_ : _06245_;
  assign _06248_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [5] : \MSYNC_1r1w.synth.nz.mem[60] [5];
  assign _06249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [5] : \MSYNC_1r1w.synth.nz.mem[62] [5];
  assign _06250_ = \bapg_rd.w_ptr_r [1] ? _06249_ : _06248_;
  assign _06251_ = \bapg_rd.w_ptr_r [2] ? _06250_ : _06247_;
  assign _06252_ = \bapg_rd.w_ptr_r [3] ? _06251_ : _06244_;
  assign _06253_ = \bapg_rd.w_ptr_r [4] ? _06252_ : _06237_;
  assign _06254_ = \bapg_rd.w_ptr_r [5] ? _06253_ : _06222_;
  assign _06255_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [5] : \MSYNC_1r1w.synth.nz.mem[64] [5];
  assign _06256_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [5] : \MSYNC_1r1w.synth.nz.mem[66] [5];
  assign _06257_ = \bapg_rd.w_ptr_r [1] ? _06256_ : _06255_;
  assign _06258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [5] : \MSYNC_1r1w.synth.nz.mem[68] [5];
  assign _06259_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [5] : \MSYNC_1r1w.synth.nz.mem[70] [5];
  assign _06260_ = \bapg_rd.w_ptr_r [1] ? _06259_ : _06258_;
  assign _06261_ = \bapg_rd.w_ptr_r [2] ? _06260_ : _06257_;
  assign _06262_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [5] : \MSYNC_1r1w.synth.nz.mem[72] [5];
  assign _06263_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [5] : \MSYNC_1r1w.synth.nz.mem[74] [5];
  assign _06264_ = \bapg_rd.w_ptr_r [1] ? _06263_ : _06262_;
  assign _06265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [5] : \MSYNC_1r1w.synth.nz.mem[76] [5];
  assign _06266_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [5] : \MSYNC_1r1w.synth.nz.mem[78] [5];
  assign _06267_ = \bapg_rd.w_ptr_r [1] ? _06266_ : _06265_;
  assign _06268_ = \bapg_rd.w_ptr_r [2] ? _06267_ : _06264_;
  assign _06269_ = \bapg_rd.w_ptr_r [3] ? _06268_ : _06261_;
  assign _06270_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [5] : \MSYNC_1r1w.synth.nz.mem[80] [5];
  assign _06271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [5] : \MSYNC_1r1w.synth.nz.mem[82] [5];
  assign _06272_ = \bapg_rd.w_ptr_r [1] ? _06271_ : _06270_;
  assign _06273_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [5] : \MSYNC_1r1w.synth.nz.mem[84] [5];
  assign _06274_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [5] : \MSYNC_1r1w.synth.nz.mem[86] [5];
  assign _06275_ = \bapg_rd.w_ptr_r [1] ? _06274_ : _06273_;
  assign _06276_ = \bapg_rd.w_ptr_r [2] ? _06275_ : _06272_;
  assign _06277_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [5] : \MSYNC_1r1w.synth.nz.mem[88] [5];
  assign _06278_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [5] : \MSYNC_1r1w.synth.nz.mem[90] [5];
  assign _06279_ = \bapg_rd.w_ptr_r [1] ? _06278_ : _06277_;
  assign _06280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [5] : \MSYNC_1r1w.synth.nz.mem[92] [5];
  assign _06281_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [5] : \MSYNC_1r1w.synth.nz.mem[94] [5];
  assign _06282_ = \bapg_rd.w_ptr_r [1] ? _06281_ : _06280_;
  assign _06283_ = \bapg_rd.w_ptr_r [2] ? _06282_ : _06279_;
  assign _06284_ = \bapg_rd.w_ptr_r [3] ? _06283_ : _06276_;
  assign _06285_ = \bapg_rd.w_ptr_r [4] ? _06284_ : _06269_;
  assign _06286_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [5] : \MSYNC_1r1w.synth.nz.mem[96] [5];
  assign _06287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [5] : \MSYNC_1r1w.synth.nz.mem[98] [5];
  assign _06288_ = \bapg_rd.w_ptr_r [1] ? _06287_ : _06286_;
  assign _06289_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [5] : \MSYNC_1r1w.synth.nz.mem[100] [5];
  assign _06290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [5] : \MSYNC_1r1w.synth.nz.mem[102] [5];
  assign _06291_ = \bapg_rd.w_ptr_r [1] ? _06290_ : _06289_;
  assign _06292_ = \bapg_rd.w_ptr_r [2] ? _06291_ : _06288_;
  assign _06293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [5] : \MSYNC_1r1w.synth.nz.mem[104] [5];
  assign _06294_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [5] : \MSYNC_1r1w.synth.nz.mem[106] [5];
  assign _06295_ = \bapg_rd.w_ptr_r [1] ? _06294_ : _06293_;
  assign _06296_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [5] : \MSYNC_1r1w.synth.nz.mem[108] [5];
  assign _06297_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [5] : \MSYNC_1r1w.synth.nz.mem[110] [5];
  assign _06298_ = \bapg_rd.w_ptr_r [1] ? _06297_ : _06296_;
  assign _06299_ = \bapg_rd.w_ptr_r [2] ? _06298_ : _06295_;
  assign _06300_ = \bapg_rd.w_ptr_r [3] ? _06299_ : _06292_;
  assign _06301_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [5] : \MSYNC_1r1w.synth.nz.mem[112] [5];
  assign _06302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [5] : \MSYNC_1r1w.synth.nz.mem[114] [5];
  assign _06303_ = \bapg_rd.w_ptr_r [1] ? _06302_ : _06301_;
  assign _06304_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [5] : \MSYNC_1r1w.synth.nz.mem[116] [5];
  assign _06305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [5] : \MSYNC_1r1w.synth.nz.mem[118] [5];
  assign _06306_ = \bapg_rd.w_ptr_r [1] ? _06305_ : _06304_;
  assign _06307_ = \bapg_rd.w_ptr_r [2] ? _06306_ : _06303_;
  assign _06308_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [5] : \MSYNC_1r1w.synth.nz.mem[120] [5];
  assign _06309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [5] : \MSYNC_1r1w.synth.nz.mem[122] [5];
  assign _06310_ = \bapg_rd.w_ptr_r [1] ? _06309_ : _06308_;
  assign _06311_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [5] : \MSYNC_1r1w.synth.nz.mem[124] [5];
  assign _06312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [5] : \MSYNC_1r1w.synth.nz.mem[126] [5];
  assign _06313_ = \bapg_rd.w_ptr_r [1] ? _06312_ : _06311_;
  assign _06314_ = \bapg_rd.w_ptr_r [2] ? _06313_ : _06310_;
  assign _06315_ = \bapg_rd.w_ptr_r [3] ? _06314_ : _06307_;
  assign _06316_ = \bapg_rd.w_ptr_r [4] ? _06315_ : _06300_;
  assign _06317_ = \bapg_rd.w_ptr_r [5] ? _06316_ : _06285_;
  assign _06318_ = \bapg_rd.w_ptr_r [6] ? _06317_ : _06254_;
  assign _06319_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [5] : \MSYNC_1r1w.synth.nz.mem[128] [5];
  assign _06320_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [5] : \MSYNC_1r1w.synth.nz.mem[130] [5];
  assign _06321_ = \bapg_rd.w_ptr_r [1] ? _06320_ : _06319_;
  assign _06322_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [5] : \MSYNC_1r1w.synth.nz.mem[132] [5];
  assign _06323_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [5] : \MSYNC_1r1w.synth.nz.mem[134] [5];
  assign _06324_ = \bapg_rd.w_ptr_r [1] ? _06323_ : _06322_;
  assign _06325_ = \bapg_rd.w_ptr_r [2] ? _06324_ : _06321_;
  assign _06326_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [5] : \MSYNC_1r1w.synth.nz.mem[136] [5];
  assign _06327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [5] : \MSYNC_1r1w.synth.nz.mem[138] [5];
  assign _06328_ = \bapg_rd.w_ptr_r [1] ? _06327_ : _06326_;
  assign _06329_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [5] : \MSYNC_1r1w.synth.nz.mem[140] [5];
  assign _06330_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [5] : \MSYNC_1r1w.synth.nz.mem[142] [5];
  assign _06331_ = \bapg_rd.w_ptr_r [1] ? _06330_ : _06329_;
  assign _06332_ = \bapg_rd.w_ptr_r [2] ? _06331_ : _06328_;
  assign _06333_ = \bapg_rd.w_ptr_r [3] ? _06332_ : _06325_;
  assign _06334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [5] : \MSYNC_1r1w.synth.nz.mem[144] [5];
  assign _06335_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [5] : \MSYNC_1r1w.synth.nz.mem[146] [5];
  assign _06336_ = \bapg_rd.w_ptr_r [1] ? _06335_ : _06334_;
  assign _06337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [5] : \MSYNC_1r1w.synth.nz.mem[148] [5];
  assign _06338_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [5] : \MSYNC_1r1w.synth.nz.mem[150] [5];
  assign _06339_ = \bapg_rd.w_ptr_r [1] ? _06338_ : _06337_;
  assign _06340_ = \bapg_rd.w_ptr_r [2] ? _06339_ : _06336_;
  assign _06341_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [5] : \MSYNC_1r1w.synth.nz.mem[152] [5];
  assign _06342_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [5] : \MSYNC_1r1w.synth.nz.mem[154] [5];
  assign _06343_ = \bapg_rd.w_ptr_r [1] ? _06342_ : _06341_;
  assign _06344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [5] : \MSYNC_1r1w.synth.nz.mem[156] [5];
  assign _06345_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [5] : \MSYNC_1r1w.synth.nz.mem[158] [5];
  assign _06346_ = \bapg_rd.w_ptr_r [1] ? _06345_ : _06344_;
  assign _06347_ = \bapg_rd.w_ptr_r [2] ? _06346_ : _06343_;
  assign _06348_ = \bapg_rd.w_ptr_r [3] ? _06347_ : _06340_;
  assign _06349_ = \bapg_rd.w_ptr_r [4] ? _06348_ : _06333_;
  assign _06350_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [5] : \MSYNC_1r1w.synth.nz.mem[160] [5];
  assign _06351_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [5] : \MSYNC_1r1w.synth.nz.mem[162] [5];
  assign _06352_ = \bapg_rd.w_ptr_r [1] ? _06351_ : _06350_;
  assign _06353_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [5] : \MSYNC_1r1w.synth.nz.mem[164] [5];
  assign _06354_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [5] : \MSYNC_1r1w.synth.nz.mem[166] [5];
  assign _06355_ = \bapg_rd.w_ptr_r [1] ? _06354_ : _06353_;
  assign _06356_ = \bapg_rd.w_ptr_r [2] ? _06355_ : _06352_;
  assign _06357_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [5] : \MSYNC_1r1w.synth.nz.mem[168] [5];
  assign _06358_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [5] : \MSYNC_1r1w.synth.nz.mem[170] [5];
  assign _06359_ = \bapg_rd.w_ptr_r [1] ? _06358_ : _06357_;
  assign _06360_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [5] : \MSYNC_1r1w.synth.nz.mem[172] [5];
  assign _06361_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [5] : \MSYNC_1r1w.synth.nz.mem[174] [5];
  assign _06362_ = \bapg_rd.w_ptr_r [1] ? _06361_ : _06360_;
  assign _06363_ = \bapg_rd.w_ptr_r [2] ? _06362_ : _06359_;
  assign _06364_ = \bapg_rd.w_ptr_r [3] ? _06363_ : _06356_;
  assign _06365_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [5] : \MSYNC_1r1w.synth.nz.mem[176] [5];
  assign _06366_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [5] : \MSYNC_1r1w.synth.nz.mem[178] [5];
  assign _06367_ = \bapg_rd.w_ptr_r [1] ? _06366_ : _06365_;
  assign _06368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [5] : \MSYNC_1r1w.synth.nz.mem[180] [5];
  assign _06369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [5] : \MSYNC_1r1w.synth.nz.mem[182] [5];
  assign _06370_ = \bapg_rd.w_ptr_r [1] ? _06369_ : _06368_;
  assign _06371_ = \bapg_rd.w_ptr_r [2] ? _06370_ : _06367_;
  assign _06372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [5] : \MSYNC_1r1w.synth.nz.mem[184] [5];
  assign _06373_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [5] : \MSYNC_1r1w.synth.nz.mem[186] [5];
  assign _06374_ = \bapg_rd.w_ptr_r [1] ? _06373_ : _06372_;
  assign _06375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [5] : \MSYNC_1r1w.synth.nz.mem[188] [5];
  assign _06376_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [5] : \MSYNC_1r1w.synth.nz.mem[190] [5];
  assign _06377_ = \bapg_rd.w_ptr_r [1] ? _06376_ : _06375_;
  assign _06378_ = \bapg_rd.w_ptr_r [2] ? _06377_ : _06374_;
  assign _06379_ = \bapg_rd.w_ptr_r [3] ? _06378_ : _06371_;
  assign _06380_ = \bapg_rd.w_ptr_r [4] ? _06379_ : _06364_;
  assign _06381_ = \bapg_rd.w_ptr_r [5] ? _06380_ : _06349_;
  assign _06382_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [5] : \MSYNC_1r1w.synth.nz.mem[192] [5];
  assign _06383_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [5] : \MSYNC_1r1w.synth.nz.mem[194] [5];
  assign _06384_ = \bapg_rd.w_ptr_r [1] ? _06383_ : _06382_;
  assign _06385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [5] : \MSYNC_1r1w.synth.nz.mem[196] [5];
  assign _06386_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [5] : \MSYNC_1r1w.synth.nz.mem[198] [5];
  assign _06387_ = \bapg_rd.w_ptr_r [1] ? _06386_ : _06385_;
  assign _06388_ = \bapg_rd.w_ptr_r [2] ? _06387_ : _06384_;
  assign _06389_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [5] : \MSYNC_1r1w.synth.nz.mem[200] [5];
  assign _06390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [5] : \MSYNC_1r1w.synth.nz.mem[202] [5];
  assign _06391_ = \bapg_rd.w_ptr_r [1] ? _06390_ : _06389_;
  assign _06392_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [5] : \MSYNC_1r1w.synth.nz.mem[204] [5];
  assign _06393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [5] : \MSYNC_1r1w.synth.nz.mem[206] [5];
  assign _06394_ = \bapg_rd.w_ptr_r [1] ? _06393_ : _06392_;
  assign _06395_ = \bapg_rd.w_ptr_r [2] ? _06394_ : _06391_;
  assign _06396_ = \bapg_rd.w_ptr_r [3] ? _06395_ : _06388_;
  assign _06397_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [5] : \MSYNC_1r1w.synth.nz.mem[208] [5];
  assign _06398_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [5] : \MSYNC_1r1w.synth.nz.mem[210] [5];
  assign _06399_ = \bapg_rd.w_ptr_r [1] ? _06398_ : _06397_;
  assign _06400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [5] : \MSYNC_1r1w.synth.nz.mem[212] [5];
  assign _06401_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [5] : \MSYNC_1r1w.synth.nz.mem[214] [5];
  assign _06402_ = \bapg_rd.w_ptr_r [1] ? _06401_ : _06400_;
  assign _06403_ = \bapg_rd.w_ptr_r [2] ? _06402_ : _06399_;
  assign _06404_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [5] : \MSYNC_1r1w.synth.nz.mem[216] [5];
  assign _06405_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [5] : \MSYNC_1r1w.synth.nz.mem[218] [5];
  assign _06406_ = \bapg_rd.w_ptr_r [1] ? _06405_ : _06404_;
  assign _06407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [5] : \MSYNC_1r1w.synth.nz.mem[220] [5];
  assign _06408_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [5] : \MSYNC_1r1w.synth.nz.mem[222] [5];
  assign _06409_ = \bapg_rd.w_ptr_r [1] ? _06408_ : _06407_;
  assign _06410_ = \bapg_rd.w_ptr_r [2] ? _06409_ : _06406_;
  assign _06411_ = \bapg_rd.w_ptr_r [3] ? _06410_ : _06403_;
  assign _06412_ = \bapg_rd.w_ptr_r [4] ? _06411_ : _06396_;
  assign _06413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [5] : \MSYNC_1r1w.synth.nz.mem[224] [5];
  assign _06414_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [5] : \MSYNC_1r1w.synth.nz.mem[226] [5];
  assign _06415_ = \bapg_rd.w_ptr_r [1] ? _06414_ : _06413_;
  assign _06416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [5] : \MSYNC_1r1w.synth.nz.mem[228] [5];
  assign _06417_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [5] : \MSYNC_1r1w.synth.nz.mem[230] [5];
  assign _06418_ = \bapg_rd.w_ptr_r [1] ? _06417_ : _06416_;
  assign _06419_ = \bapg_rd.w_ptr_r [2] ? _06418_ : _06415_;
  assign _06420_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [5] : \MSYNC_1r1w.synth.nz.mem[232] [5];
  assign _06421_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [5] : \MSYNC_1r1w.synth.nz.mem[234] [5];
  assign _06422_ = \bapg_rd.w_ptr_r [1] ? _06421_ : _06420_;
  assign _06423_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [5] : \MSYNC_1r1w.synth.nz.mem[236] [5];
  assign _06424_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [5] : \MSYNC_1r1w.synth.nz.mem[238] [5];
  assign _06425_ = \bapg_rd.w_ptr_r [1] ? _06424_ : _06423_;
  assign _06426_ = \bapg_rd.w_ptr_r [2] ? _06425_ : _06422_;
  assign _06427_ = \bapg_rd.w_ptr_r [3] ? _06426_ : _06419_;
  assign _06428_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [5] : \MSYNC_1r1w.synth.nz.mem[240] [5];
  assign _06429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [5] : \MSYNC_1r1w.synth.nz.mem[242] [5];
  assign _06430_ = \bapg_rd.w_ptr_r [1] ? _06429_ : _06428_;
  assign _06431_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [5] : \MSYNC_1r1w.synth.nz.mem[244] [5];
  assign _06432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [5] : \MSYNC_1r1w.synth.nz.mem[246] [5];
  assign _06433_ = \bapg_rd.w_ptr_r [1] ? _06432_ : _06431_;
  assign _06434_ = \bapg_rd.w_ptr_r [2] ? _06433_ : _06430_;
  assign _06435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [5] : \MSYNC_1r1w.synth.nz.mem[248] [5];
  assign _06436_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [5] : \MSYNC_1r1w.synth.nz.mem[250] [5];
  assign _06437_ = \bapg_rd.w_ptr_r [1] ? _06436_ : _06435_;
  assign _06438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [5] : \MSYNC_1r1w.synth.nz.mem[252] [5];
  assign _06439_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [5] : \MSYNC_1r1w.synth.nz.mem[254] [5];
  assign _06440_ = \bapg_rd.w_ptr_r [1] ? _06439_ : _06438_;
  assign _06441_ = \bapg_rd.w_ptr_r [2] ? _06440_ : _06437_;
  assign _06442_ = \bapg_rd.w_ptr_r [3] ? _06441_ : _06434_;
  assign _06443_ = \bapg_rd.w_ptr_r [4] ? _06442_ : _06427_;
  assign _06444_ = \bapg_rd.w_ptr_r [5] ? _06443_ : _06412_;
  assign _06445_ = \bapg_rd.w_ptr_r [6] ? _06444_ : _06381_;
  assign _06446_ = \bapg_rd.w_ptr_r [7] ? _06445_ : _06318_;
  assign _06447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [5] : \MSYNC_1r1w.synth.nz.mem[256] [5];
  assign _06448_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [5] : \MSYNC_1r1w.synth.nz.mem[258] [5];
  assign _06449_ = \bapg_rd.w_ptr_r [1] ? _06448_ : _06447_;
  assign _06450_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [5] : \MSYNC_1r1w.synth.nz.mem[260] [5];
  assign _06451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [5] : \MSYNC_1r1w.synth.nz.mem[262] [5];
  assign _06452_ = \bapg_rd.w_ptr_r [1] ? _06451_ : _06450_;
  assign _06453_ = \bapg_rd.w_ptr_r [2] ? _06452_ : _06449_;
  assign _06454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [5] : \MSYNC_1r1w.synth.nz.mem[264] [5];
  assign _06455_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [5] : \MSYNC_1r1w.synth.nz.mem[266] [5];
  assign _06456_ = \bapg_rd.w_ptr_r [1] ? _06455_ : _06454_;
  assign _06457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [5] : \MSYNC_1r1w.synth.nz.mem[268] [5];
  assign _06458_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [5] : \MSYNC_1r1w.synth.nz.mem[270] [5];
  assign _06459_ = \bapg_rd.w_ptr_r [1] ? _06458_ : _06457_;
  assign _06460_ = \bapg_rd.w_ptr_r [2] ? _06459_ : _06456_;
  assign _06461_ = \bapg_rd.w_ptr_r [3] ? _06460_ : _06453_;
  assign _06462_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [5] : \MSYNC_1r1w.synth.nz.mem[272] [5];
  assign _06463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [5] : \MSYNC_1r1w.synth.nz.mem[274] [5];
  assign _06464_ = \bapg_rd.w_ptr_r [1] ? _06463_ : _06462_;
  assign _06465_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [5] : \MSYNC_1r1w.synth.nz.mem[276] [5];
  assign _06466_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [5] : \MSYNC_1r1w.synth.nz.mem[278] [5];
  assign _06467_ = \bapg_rd.w_ptr_r [1] ? _06466_ : _06465_;
  assign _06468_ = \bapg_rd.w_ptr_r [2] ? _06467_ : _06464_;
  assign _06469_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [5] : \MSYNC_1r1w.synth.nz.mem[280] [5];
  assign _06470_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [5] : \MSYNC_1r1w.synth.nz.mem[282] [5];
  assign _06471_ = \bapg_rd.w_ptr_r [1] ? _06470_ : _06469_;
  assign _06472_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [5] : \MSYNC_1r1w.synth.nz.mem[284] [5];
  assign _06473_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [5] : \MSYNC_1r1w.synth.nz.mem[286] [5];
  assign _06474_ = \bapg_rd.w_ptr_r [1] ? _06473_ : _06472_;
  assign _06475_ = \bapg_rd.w_ptr_r [2] ? _06474_ : _06471_;
  assign _06476_ = \bapg_rd.w_ptr_r [3] ? _06475_ : _06468_;
  assign _06477_ = \bapg_rd.w_ptr_r [4] ? _06476_ : _06461_;
  assign _06478_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [5] : \MSYNC_1r1w.synth.nz.mem[288] [5];
  assign _06479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [5] : \MSYNC_1r1w.synth.nz.mem[290] [5];
  assign _06480_ = \bapg_rd.w_ptr_r [1] ? _06479_ : _06478_;
  assign _06481_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [5] : \MSYNC_1r1w.synth.nz.mem[292] [5];
  assign _06482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [5] : \MSYNC_1r1w.synth.nz.mem[294] [5];
  assign _06483_ = \bapg_rd.w_ptr_r [1] ? _06482_ : _06481_;
  assign _06484_ = \bapg_rd.w_ptr_r [2] ? _06483_ : _06480_;
  assign _06485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [5] : \MSYNC_1r1w.synth.nz.mem[296] [5];
  assign _06486_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [5] : \MSYNC_1r1w.synth.nz.mem[298] [5];
  assign _06487_ = \bapg_rd.w_ptr_r [1] ? _06486_ : _06485_;
  assign _06488_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [5] : \MSYNC_1r1w.synth.nz.mem[300] [5];
  assign _06489_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [5] : \MSYNC_1r1w.synth.nz.mem[302] [5];
  assign _06490_ = \bapg_rd.w_ptr_r [1] ? _06489_ : _06488_;
  assign _06491_ = \bapg_rd.w_ptr_r [2] ? _06490_ : _06487_;
  assign _06492_ = \bapg_rd.w_ptr_r [3] ? _06491_ : _06484_;
  assign _06493_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [5] : \MSYNC_1r1w.synth.nz.mem[304] [5];
  assign _06494_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [5] : \MSYNC_1r1w.synth.nz.mem[306] [5];
  assign _06495_ = \bapg_rd.w_ptr_r [1] ? _06494_ : _06493_;
  assign _06496_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [5] : \MSYNC_1r1w.synth.nz.mem[308] [5];
  assign _06497_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [5] : \MSYNC_1r1w.synth.nz.mem[310] [5];
  assign _06498_ = \bapg_rd.w_ptr_r [1] ? _06497_ : _06496_;
  assign _06499_ = \bapg_rd.w_ptr_r [2] ? _06498_ : _06495_;
  assign _06500_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [5] : \MSYNC_1r1w.synth.nz.mem[312] [5];
  assign _06501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [5] : \MSYNC_1r1w.synth.nz.mem[314] [5];
  assign _06502_ = \bapg_rd.w_ptr_r [1] ? _06501_ : _06500_;
  assign _06503_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [5] : \MSYNC_1r1w.synth.nz.mem[316] [5];
  assign _06504_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [5] : \MSYNC_1r1w.synth.nz.mem[318] [5];
  assign _06505_ = \bapg_rd.w_ptr_r [1] ? _06504_ : _06503_;
  assign _06506_ = \bapg_rd.w_ptr_r [2] ? _06505_ : _06502_;
  assign _06507_ = \bapg_rd.w_ptr_r [3] ? _06506_ : _06499_;
  assign _06508_ = \bapg_rd.w_ptr_r [4] ? _06507_ : _06492_;
  assign _06509_ = \bapg_rd.w_ptr_r [5] ? _06508_ : _06477_;
  assign _06510_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [5] : \MSYNC_1r1w.synth.nz.mem[320] [5];
  assign _06511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [5] : \MSYNC_1r1w.synth.nz.mem[322] [5];
  assign _06512_ = \bapg_rd.w_ptr_r [1] ? _06511_ : _06510_;
  assign _06513_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [5] : \MSYNC_1r1w.synth.nz.mem[324] [5];
  assign _06514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [5] : \MSYNC_1r1w.synth.nz.mem[326] [5];
  assign _06515_ = \bapg_rd.w_ptr_r [1] ? _06514_ : _06513_;
  assign _06516_ = \bapg_rd.w_ptr_r [2] ? _06515_ : _06512_;
  assign _06517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [5] : \MSYNC_1r1w.synth.nz.mem[328] [5];
  assign _06518_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [5] : \MSYNC_1r1w.synth.nz.mem[330] [5];
  assign _06519_ = \bapg_rd.w_ptr_r [1] ? _06518_ : _06517_;
  assign _06520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [5] : \MSYNC_1r1w.synth.nz.mem[332] [5];
  assign _06521_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [5] : \MSYNC_1r1w.synth.nz.mem[334] [5];
  assign _06522_ = \bapg_rd.w_ptr_r [1] ? _06521_ : _06520_;
  assign _06523_ = \bapg_rd.w_ptr_r [2] ? _06522_ : _06519_;
  assign _06524_ = \bapg_rd.w_ptr_r [3] ? _06523_ : _06516_;
  assign _06525_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [5] : \MSYNC_1r1w.synth.nz.mem[336] [5];
  assign _06526_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [5] : \MSYNC_1r1w.synth.nz.mem[338] [5];
  assign _06527_ = \bapg_rd.w_ptr_r [1] ? _06526_ : _06525_;
  assign _06528_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [5] : \MSYNC_1r1w.synth.nz.mem[340] [5];
  assign _06529_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [5] : \MSYNC_1r1w.synth.nz.mem[342] [5];
  assign _06530_ = \bapg_rd.w_ptr_r [1] ? _06529_ : _06528_;
  assign _06531_ = \bapg_rd.w_ptr_r [2] ? _06530_ : _06527_;
  assign _06532_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [5] : \MSYNC_1r1w.synth.nz.mem[344] [5];
  assign _06533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [5] : \MSYNC_1r1w.synth.nz.mem[346] [5];
  assign _06534_ = \bapg_rd.w_ptr_r [1] ? _06533_ : _06532_;
  assign _06535_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [5] : \MSYNC_1r1w.synth.nz.mem[348] [5];
  assign _06536_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [5] : \MSYNC_1r1w.synth.nz.mem[350] [5];
  assign _06537_ = \bapg_rd.w_ptr_r [1] ? _06536_ : _06535_;
  assign _06538_ = \bapg_rd.w_ptr_r [2] ? _06537_ : _06534_;
  assign _06539_ = \bapg_rd.w_ptr_r [3] ? _06538_ : _06531_;
  assign _06540_ = \bapg_rd.w_ptr_r [4] ? _06539_ : _06524_;
  assign _06541_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [5] : \MSYNC_1r1w.synth.nz.mem[352] [5];
  assign _06542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [5] : \MSYNC_1r1w.synth.nz.mem[354] [5];
  assign _06543_ = \bapg_rd.w_ptr_r [1] ? _06542_ : _06541_;
  assign _06544_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [5] : \MSYNC_1r1w.synth.nz.mem[356] [5];
  assign _06545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [5] : \MSYNC_1r1w.synth.nz.mem[358] [5];
  assign _06546_ = \bapg_rd.w_ptr_r [1] ? _06545_ : _06544_;
  assign _06547_ = \bapg_rd.w_ptr_r [2] ? _06546_ : _06543_;
  assign _06548_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [5] : \MSYNC_1r1w.synth.nz.mem[360] [5];
  assign _06549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [5] : \MSYNC_1r1w.synth.nz.mem[362] [5];
  assign _06550_ = \bapg_rd.w_ptr_r [1] ? _06549_ : _06548_;
  assign _06551_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [5] : \MSYNC_1r1w.synth.nz.mem[364] [5];
  assign _06552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [5] : \MSYNC_1r1w.synth.nz.mem[366] [5];
  assign _06553_ = \bapg_rd.w_ptr_r [1] ? _06552_ : _06551_;
  assign _06554_ = \bapg_rd.w_ptr_r [2] ? _06553_ : _06550_;
  assign _06555_ = \bapg_rd.w_ptr_r [3] ? _06554_ : _06547_;
  assign _06556_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [5] : \MSYNC_1r1w.synth.nz.mem[368] [5];
  assign _06557_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [5] : \MSYNC_1r1w.synth.nz.mem[370] [5];
  assign _06558_ = \bapg_rd.w_ptr_r [1] ? _06557_ : _06556_;
  assign _06559_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [5] : \MSYNC_1r1w.synth.nz.mem[372] [5];
  assign _06560_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [5] : \MSYNC_1r1w.synth.nz.mem[374] [5];
  assign _06561_ = \bapg_rd.w_ptr_r [1] ? _06560_ : _06559_;
  assign _06562_ = \bapg_rd.w_ptr_r [2] ? _06561_ : _06558_;
  assign _06563_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [5] : \MSYNC_1r1w.synth.nz.mem[376] [5];
  assign _06564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [5] : \MSYNC_1r1w.synth.nz.mem[378] [5];
  assign _06565_ = \bapg_rd.w_ptr_r [1] ? _06564_ : _06563_;
  assign _06566_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [5] : \MSYNC_1r1w.synth.nz.mem[380] [5];
  assign _06567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [5] : \MSYNC_1r1w.synth.nz.mem[382] [5];
  assign _06568_ = \bapg_rd.w_ptr_r [1] ? _06567_ : _06566_;
  assign _06569_ = \bapg_rd.w_ptr_r [2] ? _06568_ : _06565_;
  assign _06570_ = \bapg_rd.w_ptr_r [3] ? _06569_ : _06562_;
  assign _06571_ = \bapg_rd.w_ptr_r [4] ? _06570_ : _06555_;
  assign _06572_ = \bapg_rd.w_ptr_r [5] ? _06571_ : _06540_;
  assign _06573_ = \bapg_rd.w_ptr_r [6] ? _06572_ : _06509_;
  assign _06574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [5] : \MSYNC_1r1w.synth.nz.mem[384] [5];
  assign _06575_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [5] : \MSYNC_1r1w.synth.nz.mem[386] [5];
  assign _06576_ = \bapg_rd.w_ptr_r [1] ? _06575_ : _06574_;
  assign _06577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [5] : \MSYNC_1r1w.synth.nz.mem[388] [5];
  assign _06578_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [5] : \MSYNC_1r1w.synth.nz.mem[390] [5];
  assign _06579_ = \bapg_rd.w_ptr_r [1] ? _06578_ : _06577_;
  assign _06580_ = \bapg_rd.w_ptr_r [2] ? _06579_ : _06576_;
  assign _06581_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [5] : \MSYNC_1r1w.synth.nz.mem[392] [5];
  assign _06582_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [5] : \MSYNC_1r1w.synth.nz.mem[394] [5];
  assign _06583_ = \bapg_rd.w_ptr_r [1] ? _06582_ : _06581_;
  assign _06584_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [5] : \MSYNC_1r1w.synth.nz.mem[396] [5];
  assign _06585_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [5] : \MSYNC_1r1w.synth.nz.mem[398] [5];
  assign _06586_ = \bapg_rd.w_ptr_r [1] ? _06585_ : _06584_;
  assign _06587_ = \bapg_rd.w_ptr_r [2] ? _06586_ : _06583_;
  assign _06588_ = \bapg_rd.w_ptr_r [3] ? _06587_ : _06580_;
  assign _06589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [5] : \MSYNC_1r1w.synth.nz.mem[400] [5];
  assign _06590_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [5] : \MSYNC_1r1w.synth.nz.mem[402] [5];
  assign _06591_ = \bapg_rd.w_ptr_r [1] ? _06590_ : _06589_;
  assign _06592_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [5] : \MSYNC_1r1w.synth.nz.mem[404] [5];
  assign _06593_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [5] : \MSYNC_1r1w.synth.nz.mem[406] [5];
  assign _06594_ = \bapg_rd.w_ptr_r [1] ? _06593_ : _06592_;
  assign _06595_ = \bapg_rd.w_ptr_r [2] ? _06594_ : _06591_;
  assign _06596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [5] : \MSYNC_1r1w.synth.nz.mem[408] [5];
  assign _06597_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [5] : \MSYNC_1r1w.synth.nz.mem[410] [5];
  assign _06598_ = \bapg_rd.w_ptr_r [1] ? _06597_ : _06596_;
  assign _06599_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [5] : \MSYNC_1r1w.synth.nz.mem[412] [5];
  assign _06600_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [5] : \MSYNC_1r1w.synth.nz.mem[414] [5];
  assign _06601_ = \bapg_rd.w_ptr_r [1] ? _06600_ : _06599_;
  assign _06602_ = \bapg_rd.w_ptr_r [2] ? _06601_ : _06598_;
  assign _06603_ = \bapg_rd.w_ptr_r [3] ? _06602_ : _06595_;
  assign _06604_ = \bapg_rd.w_ptr_r [4] ? _06603_ : _06588_;
  assign _06605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [5] : \MSYNC_1r1w.synth.nz.mem[416] [5];
  assign _06606_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [5] : \MSYNC_1r1w.synth.nz.mem[418] [5];
  assign _06607_ = \bapg_rd.w_ptr_r [1] ? _06606_ : _06605_;
  assign _06608_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [5] : \MSYNC_1r1w.synth.nz.mem[420] [5];
  assign _06609_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [5] : \MSYNC_1r1w.synth.nz.mem[422] [5];
  assign _06610_ = \bapg_rd.w_ptr_r [1] ? _06609_ : _06608_;
  assign _06611_ = \bapg_rd.w_ptr_r [2] ? _06610_ : _06607_;
  assign _06612_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [5] : \MSYNC_1r1w.synth.nz.mem[424] [5];
  assign _06613_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [5] : \MSYNC_1r1w.synth.nz.mem[426] [5];
  assign _06614_ = \bapg_rd.w_ptr_r [1] ? _06613_ : _06612_;
  assign _06615_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [5] : \MSYNC_1r1w.synth.nz.mem[428] [5];
  assign _06616_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [5] : \MSYNC_1r1w.synth.nz.mem[430] [5];
  assign _06617_ = \bapg_rd.w_ptr_r [1] ? _06616_ : _06615_;
  assign _06618_ = \bapg_rd.w_ptr_r [2] ? _06617_ : _06614_;
  assign _06619_ = \bapg_rd.w_ptr_r [3] ? _06618_ : _06611_;
  assign _06620_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [5] : \MSYNC_1r1w.synth.nz.mem[432] [5];
  assign _06621_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [5] : \MSYNC_1r1w.synth.nz.mem[434] [5];
  assign _06622_ = \bapg_rd.w_ptr_r [1] ? _06621_ : _06620_;
  assign _06623_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [5] : \MSYNC_1r1w.synth.nz.mem[436] [5];
  assign _06624_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [5] : \MSYNC_1r1w.synth.nz.mem[438] [5];
  assign _06625_ = \bapg_rd.w_ptr_r [1] ? _06624_ : _06623_;
  assign _06626_ = \bapg_rd.w_ptr_r [2] ? _06625_ : _06622_;
  assign _06627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [5] : \MSYNC_1r1w.synth.nz.mem[440] [5];
  assign _06628_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [5] : \MSYNC_1r1w.synth.nz.mem[442] [5];
  assign _06629_ = \bapg_rd.w_ptr_r [1] ? _06628_ : _06627_;
  assign _06630_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [5] : \MSYNC_1r1w.synth.nz.mem[444] [5];
  assign _06631_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [5] : \MSYNC_1r1w.synth.nz.mem[446] [5];
  assign _06632_ = \bapg_rd.w_ptr_r [1] ? _06631_ : _06630_;
  assign _06633_ = \bapg_rd.w_ptr_r [2] ? _06632_ : _06629_;
  assign _06634_ = \bapg_rd.w_ptr_r [3] ? _06633_ : _06626_;
  assign _06635_ = \bapg_rd.w_ptr_r [4] ? _06634_ : _06619_;
  assign _06636_ = \bapg_rd.w_ptr_r [5] ? _06635_ : _06604_;
  assign _06637_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [5] : \MSYNC_1r1w.synth.nz.mem[448] [5];
  assign _06638_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [5] : \MSYNC_1r1w.synth.nz.mem[450] [5];
  assign _06639_ = \bapg_rd.w_ptr_r [1] ? _06638_ : _06637_;
  assign _06640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [5] : \MSYNC_1r1w.synth.nz.mem[452] [5];
  assign _06641_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [5] : \MSYNC_1r1w.synth.nz.mem[454] [5];
  assign _06642_ = \bapg_rd.w_ptr_r [1] ? _06641_ : _06640_;
  assign _06643_ = \bapg_rd.w_ptr_r [2] ? _06642_ : _06639_;
  assign _06644_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [5] : \MSYNC_1r1w.synth.nz.mem[456] [5];
  assign _06645_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [5] : \MSYNC_1r1w.synth.nz.mem[458] [5];
  assign _06646_ = \bapg_rd.w_ptr_r [1] ? _06645_ : _06644_;
  assign _06647_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [5] : \MSYNC_1r1w.synth.nz.mem[460] [5];
  assign _06648_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [5] : \MSYNC_1r1w.synth.nz.mem[462] [5];
  assign _06649_ = \bapg_rd.w_ptr_r [1] ? _06648_ : _06647_;
  assign _06650_ = \bapg_rd.w_ptr_r [2] ? _06649_ : _06646_;
  assign _06651_ = \bapg_rd.w_ptr_r [3] ? _06650_ : _06643_;
  assign _06652_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [5] : \MSYNC_1r1w.synth.nz.mem[464] [5];
  assign _06653_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [5] : \MSYNC_1r1w.synth.nz.mem[466] [5];
  assign _06654_ = \bapg_rd.w_ptr_r [1] ? _06653_ : _06652_;
  assign _06655_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [5] : \MSYNC_1r1w.synth.nz.mem[468] [5];
  assign _06656_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [5] : \MSYNC_1r1w.synth.nz.mem[470] [5];
  assign _06657_ = \bapg_rd.w_ptr_r [1] ? _06656_ : _06655_;
  assign _06658_ = \bapg_rd.w_ptr_r [2] ? _06657_ : _06654_;
  assign _06659_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [5] : \MSYNC_1r1w.synth.nz.mem[472] [5];
  assign _06660_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [5] : \MSYNC_1r1w.synth.nz.mem[474] [5];
  assign _06661_ = \bapg_rd.w_ptr_r [1] ? _06660_ : _06659_;
  assign _06662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [5] : \MSYNC_1r1w.synth.nz.mem[476] [5];
  assign _06663_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [5] : \MSYNC_1r1w.synth.nz.mem[478] [5];
  assign _06664_ = \bapg_rd.w_ptr_r [1] ? _06663_ : _06662_;
  assign _06665_ = \bapg_rd.w_ptr_r [2] ? _06664_ : _06661_;
  assign _06666_ = \bapg_rd.w_ptr_r [3] ? _06665_ : _06658_;
  assign _06667_ = \bapg_rd.w_ptr_r [4] ? _06666_ : _06651_;
  assign _06668_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [5] : \MSYNC_1r1w.synth.nz.mem[480] [5];
  assign _06669_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [5] : \MSYNC_1r1w.synth.nz.mem[482] [5];
  assign _06670_ = \bapg_rd.w_ptr_r [1] ? _06669_ : _06668_;
  assign _06671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [5] : \MSYNC_1r1w.synth.nz.mem[484] [5];
  assign _06672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [5] : \MSYNC_1r1w.synth.nz.mem[486] [5];
  assign _06673_ = \bapg_rd.w_ptr_r [1] ? _06672_ : _06671_;
  assign _06674_ = \bapg_rd.w_ptr_r [2] ? _06673_ : _06670_;
  assign _06675_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [5] : \MSYNC_1r1w.synth.nz.mem[488] [5];
  assign _06676_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [5] : \MSYNC_1r1w.synth.nz.mem[490] [5];
  assign _06677_ = \bapg_rd.w_ptr_r [1] ? _06676_ : _06675_;
  assign _06678_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [5] : \MSYNC_1r1w.synth.nz.mem[492] [5];
  assign _06679_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [5] : \MSYNC_1r1w.synth.nz.mem[494] [5];
  assign _06680_ = \bapg_rd.w_ptr_r [1] ? _06679_ : _06678_;
  assign _06681_ = \bapg_rd.w_ptr_r [2] ? _06680_ : _06677_;
  assign _06682_ = \bapg_rd.w_ptr_r [3] ? _06681_ : _06674_;
  assign _06683_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [5] : \MSYNC_1r1w.synth.nz.mem[496] [5];
  assign _06684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [5] : \MSYNC_1r1w.synth.nz.mem[498] [5];
  assign _06685_ = \bapg_rd.w_ptr_r [1] ? _06684_ : _06683_;
  assign _06686_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [5] : \MSYNC_1r1w.synth.nz.mem[500] [5];
  assign _06687_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [5] : \MSYNC_1r1w.synth.nz.mem[502] [5];
  assign _06688_ = \bapg_rd.w_ptr_r [1] ? _06687_ : _06686_;
  assign _06689_ = \bapg_rd.w_ptr_r [2] ? _06688_ : _06685_;
  assign _06690_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [5] : \MSYNC_1r1w.synth.nz.mem[504] [5];
  assign _06691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [5] : \MSYNC_1r1w.synth.nz.mem[506] [5];
  assign _06692_ = \bapg_rd.w_ptr_r [1] ? _06691_ : _06690_;
  assign _06693_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [5] : \MSYNC_1r1w.synth.nz.mem[508] [5];
  assign _06694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [5] : \MSYNC_1r1w.synth.nz.mem[510] [5];
  assign _06695_ = \bapg_rd.w_ptr_r [1] ? _06694_ : _06693_;
  assign _06696_ = \bapg_rd.w_ptr_r [2] ? _06695_ : _06692_;
  assign _06697_ = \bapg_rd.w_ptr_r [3] ? _06696_ : _06689_;
  assign _06698_ = \bapg_rd.w_ptr_r [4] ? _06697_ : _06682_;
  assign _06699_ = \bapg_rd.w_ptr_r [5] ? _06698_ : _06667_;
  assign _06700_ = \bapg_rd.w_ptr_r [6] ? _06699_ : _06636_;
  assign _06701_ = \bapg_rd.w_ptr_r [7] ? _06700_ : _06573_;
  assign _06702_ = \bapg_rd.w_ptr_r [8] ? _06701_ : _06446_;
  assign _06703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [5] : \MSYNC_1r1w.synth.nz.mem[512] [5];
  assign _06704_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [5] : \MSYNC_1r1w.synth.nz.mem[514] [5];
  assign _06705_ = \bapg_rd.w_ptr_r [1] ? _06704_ : _06703_;
  assign _06706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [5] : \MSYNC_1r1w.synth.nz.mem[516] [5];
  assign _06707_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [5] : \MSYNC_1r1w.synth.nz.mem[518] [5];
  assign _06708_ = \bapg_rd.w_ptr_r [1] ? _06707_ : _06706_;
  assign _06709_ = \bapg_rd.w_ptr_r [2] ? _06708_ : _06705_;
  assign _06710_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [5] : \MSYNC_1r1w.synth.nz.mem[520] [5];
  assign _06711_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [5] : \MSYNC_1r1w.synth.nz.mem[522] [5];
  assign _06712_ = \bapg_rd.w_ptr_r [1] ? _06711_ : _06710_;
  assign _06713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [5] : \MSYNC_1r1w.synth.nz.mem[524] [5];
  assign _06714_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [5] : \MSYNC_1r1w.synth.nz.mem[526] [5];
  assign _06715_ = \bapg_rd.w_ptr_r [1] ? _06714_ : _06713_;
  assign _06716_ = \bapg_rd.w_ptr_r [2] ? _06715_ : _06712_;
  assign _06717_ = \bapg_rd.w_ptr_r [3] ? _06716_ : _06709_;
  assign _06718_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [5] : \MSYNC_1r1w.synth.nz.mem[528] [5];
  assign _06719_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [5] : \MSYNC_1r1w.synth.nz.mem[530] [5];
  assign _06720_ = \bapg_rd.w_ptr_r [1] ? _06719_ : _06718_;
  assign _06721_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [5] : \MSYNC_1r1w.synth.nz.mem[532] [5];
  assign _06722_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [5] : \MSYNC_1r1w.synth.nz.mem[534] [5];
  assign _06723_ = \bapg_rd.w_ptr_r [1] ? _06722_ : _06721_;
  assign _06724_ = \bapg_rd.w_ptr_r [2] ? _06723_ : _06720_;
  assign _06725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [5] : \MSYNC_1r1w.synth.nz.mem[536] [5];
  assign _06726_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [5] : \MSYNC_1r1w.synth.nz.mem[538] [5];
  assign _06727_ = \bapg_rd.w_ptr_r [1] ? _06726_ : _06725_;
  assign _06728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [5] : \MSYNC_1r1w.synth.nz.mem[540] [5];
  assign _06729_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [5] : \MSYNC_1r1w.synth.nz.mem[542] [5];
  assign _06730_ = \bapg_rd.w_ptr_r [1] ? _06729_ : _06728_;
  assign _06731_ = \bapg_rd.w_ptr_r [2] ? _06730_ : _06727_;
  assign _06732_ = \bapg_rd.w_ptr_r [3] ? _06731_ : _06724_;
  assign _06733_ = \bapg_rd.w_ptr_r [4] ? _06732_ : _06717_;
  assign _06734_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [5] : \MSYNC_1r1w.synth.nz.mem[544] [5];
  assign _06735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [5] : \MSYNC_1r1w.synth.nz.mem[546] [5];
  assign _06736_ = \bapg_rd.w_ptr_r [1] ? _06735_ : _06734_;
  assign _06737_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [5] : \MSYNC_1r1w.synth.nz.mem[548] [5];
  assign _06738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [5] : \MSYNC_1r1w.synth.nz.mem[550] [5];
  assign _06739_ = \bapg_rd.w_ptr_r [1] ? _06738_ : _06737_;
  assign _06740_ = \bapg_rd.w_ptr_r [2] ? _06739_ : _06736_;
  assign _06741_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [5] : \MSYNC_1r1w.synth.nz.mem[552] [5];
  assign _06742_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [5] : \MSYNC_1r1w.synth.nz.mem[554] [5];
  assign _06743_ = \bapg_rd.w_ptr_r [1] ? _06742_ : _06741_;
  assign _06744_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [5] : \MSYNC_1r1w.synth.nz.mem[556] [5];
  assign _06745_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [5] : \MSYNC_1r1w.synth.nz.mem[558] [5];
  assign _06746_ = \bapg_rd.w_ptr_r [1] ? _06745_ : _06744_;
  assign _06747_ = \bapg_rd.w_ptr_r [2] ? _06746_ : _06743_;
  assign _06748_ = \bapg_rd.w_ptr_r [3] ? _06747_ : _06740_;
  assign _06749_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [5] : \MSYNC_1r1w.synth.nz.mem[560] [5];
  assign _06750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [5] : \MSYNC_1r1w.synth.nz.mem[562] [5];
  assign _06751_ = \bapg_rd.w_ptr_r [1] ? _06750_ : _06749_;
  assign _06752_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [5] : \MSYNC_1r1w.synth.nz.mem[564] [5];
  assign _06753_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [5] : \MSYNC_1r1w.synth.nz.mem[566] [5];
  assign _06754_ = \bapg_rd.w_ptr_r [1] ? _06753_ : _06752_;
  assign _06755_ = \bapg_rd.w_ptr_r [2] ? _06754_ : _06751_;
  assign _06756_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [5] : \MSYNC_1r1w.synth.nz.mem[568] [5];
  assign _06757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [5] : \MSYNC_1r1w.synth.nz.mem[570] [5];
  assign _06758_ = \bapg_rd.w_ptr_r [1] ? _06757_ : _06756_;
  assign _06759_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [5] : \MSYNC_1r1w.synth.nz.mem[572] [5];
  assign _06760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [5] : \MSYNC_1r1w.synth.nz.mem[574] [5];
  assign _06761_ = \bapg_rd.w_ptr_r [1] ? _06760_ : _06759_;
  assign _06762_ = \bapg_rd.w_ptr_r [2] ? _06761_ : _06758_;
  assign _06763_ = \bapg_rd.w_ptr_r [3] ? _06762_ : _06755_;
  assign _06764_ = \bapg_rd.w_ptr_r [4] ? _06763_ : _06748_;
  assign _06765_ = \bapg_rd.w_ptr_r [5] ? _06764_ : _06733_;
  assign _06766_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [5] : \MSYNC_1r1w.synth.nz.mem[576] [5];
  assign _06767_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [5] : \MSYNC_1r1w.synth.nz.mem[578] [5];
  assign _06768_ = \bapg_rd.w_ptr_r [1] ? _06767_ : _06766_;
  assign _06769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [5] : \MSYNC_1r1w.synth.nz.mem[580] [5];
  assign _06770_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [5] : \MSYNC_1r1w.synth.nz.mem[582] [5];
  assign _06771_ = \bapg_rd.w_ptr_r [1] ? _06770_ : _06769_;
  assign _06772_ = \bapg_rd.w_ptr_r [2] ? _06771_ : _06768_;
  assign _06773_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [5] : \MSYNC_1r1w.synth.nz.mem[584] [5];
  assign _06774_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [5] : \MSYNC_1r1w.synth.nz.mem[586] [5];
  assign _06775_ = \bapg_rd.w_ptr_r [1] ? _06774_ : _06773_;
  assign _06776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [5] : \MSYNC_1r1w.synth.nz.mem[588] [5];
  assign _06777_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [5] : \MSYNC_1r1w.synth.nz.mem[590] [5];
  assign _06778_ = \bapg_rd.w_ptr_r [1] ? _06777_ : _06776_;
  assign _06779_ = \bapg_rd.w_ptr_r [2] ? _06778_ : _06775_;
  assign _06780_ = \bapg_rd.w_ptr_r [3] ? _06779_ : _06772_;
  assign _06781_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [5] : \MSYNC_1r1w.synth.nz.mem[592] [5];
  assign _06782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [5] : \MSYNC_1r1w.synth.nz.mem[594] [5];
  assign _06783_ = \bapg_rd.w_ptr_r [1] ? _06782_ : _06781_;
  assign _06784_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [5] : \MSYNC_1r1w.synth.nz.mem[596] [5];
  assign _06785_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [5] : \MSYNC_1r1w.synth.nz.mem[598] [5];
  assign _06786_ = \bapg_rd.w_ptr_r [1] ? _06785_ : _06784_;
  assign _06787_ = \bapg_rd.w_ptr_r [2] ? _06786_ : _06783_;
  assign _06788_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [5] : \MSYNC_1r1w.synth.nz.mem[600] [5];
  assign _06789_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [5] : \MSYNC_1r1w.synth.nz.mem[602] [5];
  assign _06790_ = \bapg_rd.w_ptr_r [1] ? _06789_ : _06788_;
  assign _06791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [5] : \MSYNC_1r1w.synth.nz.mem[604] [5];
  assign _06792_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [5] : \MSYNC_1r1w.synth.nz.mem[606] [5];
  assign _06793_ = \bapg_rd.w_ptr_r [1] ? _06792_ : _06791_;
  assign _06794_ = \bapg_rd.w_ptr_r [2] ? _06793_ : _06790_;
  assign _06795_ = \bapg_rd.w_ptr_r [3] ? _06794_ : _06787_;
  assign _06796_ = \bapg_rd.w_ptr_r [4] ? _06795_ : _06780_;
  assign _06797_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [5] : \MSYNC_1r1w.synth.nz.mem[608] [5];
  assign _06798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [5] : \MSYNC_1r1w.synth.nz.mem[610] [5];
  assign _06799_ = \bapg_rd.w_ptr_r [1] ? _06798_ : _06797_;
  assign _06800_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [5] : \MSYNC_1r1w.synth.nz.mem[612] [5];
  assign _06801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [5] : \MSYNC_1r1w.synth.nz.mem[614] [5];
  assign _06802_ = \bapg_rd.w_ptr_r [1] ? _06801_ : _06800_;
  assign _06803_ = \bapg_rd.w_ptr_r [2] ? _06802_ : _06799_;
  assign _06804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [5] : \MSYNC_1r1w.synth.nz.mem[616] [5];
  assign _06805_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [5] : \MSYNC_1r1w.synth.nz.mem[618] [5];
  assign _06806_ = \bapg_rd.w_ptr_r [1] ? _06805_ : _06804_;
  assign _06807_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [5] : \MSYNC_1r1w.synth.nz.mem[620] [5];
  assign _06808_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [5] : \MSYNC_1r1w.synth.nz.mem[622] [5];
  assign _06809_ = \bapg_rd.w_ptr_r [1] ? _06808_ : _06807_;
  assign _06810_ = \bapg_rd.w_ptr_r [2] ? _06809_ : _06806_;
  assign _06811_ = \bapg_rd.w_ptr_r [3] ? _06810_ : _06803_;
  assign _06812_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [5] : \MSYNC_1r1w.synth.nz.mem[624] [5];
  assign _06813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [5] : \MSYNC_1r1w.synth.nz.mem[626] [5];
  assign _06814_ = \bapg_rd.w_ptr_r [1] ? _06813_ : _06812_;
  assign _06815_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [5] : \MSYNC_1r1w.synth.nz.mem[628] [5];
  assign _06816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [5] : \MSYNC_1r1w.synth.nz.mem[630] [5];
  assign _06817_ = \bapg_rd.w_ptr_r [1] ? _06816_ : _06815_;
  assign _06818_ = \bapg_rd.w_ptr_r [2] ? _06817_ : _06814_;
  assign _06819_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [5] : \MSYNC_1r1w.synth.nz.mem[632] [5];
  assign _06820_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [5] : \MSYNC_1r1w.synth.nz.mem[634] [5];
  assign _06821_ = \bapg_rd.w_ptr_r [1] ? _06820_ : _06819_;
  assign _06822_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [5] : \MSYNC_1r1w.synth.nz.mem[636] [5];
  assign _06823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [5] : \MSYNC_1r1w.synth.nz.mem[638] [5];
  assign _06824_ = \bapg_rd.w_ptr_r [1] ? _06823_ : _06822_;
  assign _06825_ = \bapg_rd.w_ptr_r [2] ? _06824_ : _06821_;
  assign _06826_ = \bapg_rd.w_ptr_r [3] ? _06825_ : _06818_;
  assign _06827_ = \bapg_rd.w_ptr_r [4] ? _06826_ : _06811_;
  assign _06828_ = \bapg_rd.w_ptr_r [5] ? _06827_ : _06796_;
  assign _06829_ = \bapg_rd.w_ptr_r [6] ? _06828_ : _06765_;
  assign _06830_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [5] : \MSYNC_1r1w.synth.nz.mem[640] [5];
  assign _06831_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [5] : \MSYNC_1r1w.synth.nz.mem[642] [5];
  assign _06832_ = \bapg_rd.w_ptr_r [1] ? _06831_ : _06830_;
  assign _06833_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [5] : \MSYNC_1r1w.synth.nz.mem[644] [5];
  assign _06834_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [5] : \MSYNC_1r1w.synth.nz.mem[646] [5];
  assign _06835_ = \bapg_rd.w_ptr_r [1] ? _06834_ : _06833_;
  assign _06836_ = \bapg_rd.w_ptr_r [2] ? _06835_ : _06832_;
  assign _06837_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [5] : \MSYNC_1r1w.synth.nz.mem[648] [5];
  assign _06838_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [5] : \MSYNC_1r1w.synth.nz.mem[650] [5];
  assign _06839_ = \bapg_rd.w_ptr_r [1] ? _06838_ : _06837_;
  assign _06840_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [5] : \MSYNC_1r1w.synth.nz.mem[652] [5];
  assign _06841_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [5] : \MSYNC_1r1w.synth.nz.mem[654] [5];
  assign _06842_ = \bapg_rd.w_ptr_r [1] ? _06841_ : _06840_;
  assign _06843_ = \bapg_rd.w_ptr_r [2] ? _06842_ : _06839_;
  assign _06844_ = \bapg_rd.w_ptr_r [3] ? _06843_ : _06836_;
  assign _06845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [5] : \MSYNC_1r1w.synth.nz.mem[656] [5];
  assign _06846_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [5] : \MSYNC_1r1w.synth.nz.mem[658] [5];
  assign _06847_ = \bapg_rd.w_ptr_r [1] ? _06846_ : _06845_;
  assign _06848_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [5] : \MSYNC_1r1w.synth.nz.mem[660] [5];
  assign _06849_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [5] : \MSYNC_1r1w.synth.nz.mem[662] [5];
  assign _06850_ = \bapg_rd.w_ptr_r [1] ? _06849_ : _06848_;
  assign _06851_ = \bapg_rd.w_ptr_r [2] ? _06850_ : _06847_;
  assign _06852_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [5] : \MSYNC_1r1w.synth.nz.mem[664] [5];
  assign _06853_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [5] : \MSYNC_1r1w.synth.nz.mem[666] [5];
  assign _06854_ = \bapg_rd.w_ptr_r [1] ? _06853_ : _06852_;
  assign _06855_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [5] : \MSYNC_1r1w.synth.nz.mem[668] [5];
  assign _06856_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [5] : \MSYNC_1r1w.synth.nz.mem[670] [5];
  assign _06857_ = \bapg_rd.w_ptr_r [1] ? _06856_ : _06855_;
  assign _06858_ = \bapg_rd.w_ptr_r [2] ? _06857_ : _06854_;
  assign _06859_ = \bapg_rd.w_ptr_r [3] ? _06858_ : _06851_;
  assign _06860_ = \bapg_rd.w_ptr_r [4] ? _06859_ : _06844_;
  assign _06861_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [5] : \MSYNC_1r1w.synth.nz.mem[672] [5];
  assign _06862_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [5] : \MSYNC_1r1w.synth.nz.mem[674] [5];
  assign _06863_ = \bapg_rd.w_ptr_r [1] ? _06862_ : _06861_;
  assign _06864_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [5] : \MSYNC_1r1w.synth.nz.mem[676] [5];
  assign _06865_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [5] : \MSYNC_1r1w.synth.nz.mem[678] [5];
  assign _06866_ = \bapg_rd.w_ptr_r [1] ? _06865_ : _06864_;
  assign _06867_ = \bapg_rd.w_ptr_r [2] ? _06866_ : _06863_;
  assign _06868_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [5] : \MSYNC_1r1w.synth.nz.mem[680] [5];
  assign _06869_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [5] : \MSYNC_1r1w.synth.nz.mem[682] [5];
  assign _06870_ = \bapg_rd.w_ptr_r [1] ? _06869_ : _06868_;
  assign _06871_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [5] : \MSYNC_1r1w.synth.nz.mem[684] [5];
  assign _06872_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [5] : \MSYNC_1r1w.synth.nz.mem[686] [5];
  assign _06873_ = \bapg_rd.w_ptr_r [1] ? _06872_ : _06871_;
  assign _06874_ = \bapg_rd.w_ptr_r [2] ? _06873_ : _06870_;
  assign _06875_ = \bapg_rd.w_ptr_r [3] ? _06874_ : _06867_;
  assign _06876_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [5] : \MSYNC_1r1w.synth.nz.mem[688] [5];
  assign _06877_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [5] : \MSYNC_1r1w.synth.nz.mem[690] [5];
  assign _06878_ = \bapg_rd.w_ptr_r [1] ? _06877_ : _06876_;
  assign _06879_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [5] : \MSYNC_1r1w.synth.nz.mem[692] [5];
  assign _06880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [5] : \MSYNC_1r1w.synth.nz.mem[694] [5];
  assign _06881_ = \bapg_rd.w_ptr_r [1] ? _06880_ : _06879_;
  assign _06882_ = \bapg_rd.w_ptr_r [2] ? _06881_ : _06878_;
  assign _06883_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [5] : \MSYNC_1r1w.synth.nz.mem[696] [5];
  assign _06884_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [5] : \MSYNC_1r1w.synth.nz.mem[698] [5];
  assign _06885_ = \bapg_rd.w_ptr_r [1] ? _06884_ : _06883_;
  assign _06886_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [5] : \MSYNC_1r1w.synth.nz.mem[700] [5];
  assign _06887_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [5] : \MSYNC_1r1w.synth.nz.mem[702] [5];
  assign _06888_ = \bapg_rd.w_ptr_r [1] ? _06887_ : _06886_;
  assign _06889_ = \bapg_rd.w_ptr_r [2] ? _06888_ : _06885_;
  assign _06890_ = \bapg_rd.w_ptr_r [3] ? _06889_ : _06882_;
  assign _06891_ = \bapg_rd.w_ptr_r [4] ? _06890_ : _06875_;
  assign _06892_ = \bapg_rd.w_ptr_r [5] ? _06891_ : _06860_;
  assign _06893_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [5] : \MSYNC_1r1w.synth.nz.mem[704] [5];
  assign _06894_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [5] : \MSYNC_1r1w.synth.nz.mem[706] [5];
  assign _06895_ = \bapg_rd.w_ptr_r [1] ? _06894_ : _06893_;
  assign _06896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [5] : \MSYNC_1r1w.synth.nz.mem[708] [5];
  assign _06897_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [5] : \MSYNC_1r1w.synth.nz.mem[710] [5];
  assign _06898_ = \bapg_rd.w_ptr_r [1] ? _06897_ : _06896_;
  assign _06899_ = \bapg_rd.w_ptr_r [2] ? _06898_ : _06895_;
  assign _06900_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [5] : \MSYNC_1r1w.synth.nz.mem[712] [5];
  assign _06901_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [5] : \MSYNC_1r1w.synth.nz.mem[714] [5];
  assign _06902_ = \bapg_rd.w_ptr_r [1] ? _06901_ : _06900_;
  assign _06903_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [5] : \MSYNC_1r1w.synth.nz.mem[716] [5];
  assign _06904_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [5] : \MSYNC_1r1w.synth.nz.mem[718] [5];
  assign _06905_ = \bapg_rd.w_ptr_r [1] ? _06904_ : _06903_;
  assign _06906_ = \bapg_rd.w_ptr_r [2] ? _06905_ : _06902_;
  assign _06907_ = \bapg_rd.w_ptr_r [3] ? _06906_ : _06899_;
  assign _06908_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [5] : \MSYNC_1r1w.synth.nz.mem[720] [5];
  assign _06909_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [5] : \MSYNC_1r1w.synth.nz.mem[722] [5];
  assign _06910_ = \bapg_rd.w_ptr_r [1] ? _06909_ : _06908_;
  assign _06911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [5] : \MSYNC_1r1w.synth.nz.mem[724] [5];
  assign _06912_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [5] : \MSYNC_1r1w.synth.nz.mem[726] [5];
  assign _06913_ = \bapg_rd.w_ptr_r [1] ? _06912_ : _06911_;
  assign _06914_ = \bapg_rd.w_ptr_r [2] ? _06913_ : _06910_;
  assign _06915_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [5] : \MSYNC_1r1w.synth.nz.mem[728] [5];
  assign _06916_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [5] : \MSYNC_1r1w.synth.nz.mem[730] [5];
  assign _06917_ = \bapg_rd.w_ptr_r [1] ? _06916_ : _06915_;
  assign _06918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [5] : \MSYNC_1r1w.synth.nz.mem[732] [5];
  assign _06919_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [5] : \MSYNC_1r1w.synth.nz.mem[734] [5];
  assign _06920_ = \bapg_rd.w_ptr_r [1] ? _06919_ : _06918_;
  assign _06921_ = \bapg_rd.w_ptr_r [2] ? _06920_ : _06917_;
  assign _06922_ = \bapg_rd.w_ptr_r [3] ? _06921_ : _06914_;
  assign _06923_ = \bapg_rd.w_ptr_r [4] ? _06922_ : _06907_;
  assign _06924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [5] : \MSYNC_1r1w.synth.nz.mem[736] [5];
  assign _06925_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [5] : \MSYNC_1r1w.synth.nz.mem[738] [5];
  assign _06926_ = \bapg_rd.w_ptr_r [1] ? _06925_ : _06924_;
  assign _06927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [5] : \MSYNC_1r1w.synth.nz.mem[740] [5];
  assign _06928_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [5] : \MSYNC_1r1w.synth.nz.mem[742] [5];
  assign _06929_ = \bapg_rd.w_ptr_r [1] ? _06928_ : _06927_;
  assign _06930_ = \bapg_rd.w_ptr_r [2] ? _06929_ : _06926_;
  assign _06931_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [5] : \MSYNC_1r1w.synth.nz.mem[744] [5];
  assign _06932_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [5] : \MSYNC_1r1w.synth.nz.mem[746] [5];
  assign _06933_ = \bapg_rd.w_ptr_r [1] ? _06932_ : _06931_;
  assign _06934_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [5] : \MSYNC_1r1w.synth.nz.mem[748] [5];
  assign _06935_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [5] : \MSYNC_1r1w.synth.nz.mem[750] [5];
  assign _06936_ = \bapg_rd.w_ptr_r [1] ? _06935_ : _06934_;
  assign _06937_ = \bapg_rd.w_ptr_r [2] ? _06936_ : _06933_;
  assign _06938_ = \bapg_rd.w_ptr_r [3] ? _06937_ : _06930_;
  assign _06939_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [5] : \MSYNC_1r1w.synth.nz.mem[752] [5];
  assign _06940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [5] : \MSYNC_1r1w.synth.nz.mem[754] [5];
  assign _06941_ = \bapg_rd.w_ptr_r [1] ? _06940_ : _06939_;
  assign _06942_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [5] : \MSYNC_1r1w.synth.nz.mem[756] [5];
  assign _06943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [5] : \MSYNC_1r1w.synth.nz.mem[758] [5];
  assign _06944_ = \bapg_rd.w_ptr_r [1] ? _06943_ : _06942_;
  assign _06945_ = \bapg_rd.w_ptr_r [2] ? _06944_ : _06941_;
  assign _06946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [5] : \MSYNC_1r1w.synth.nz.mem[760] [5];
  assign _06947_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [5] : \MSYNC_1r1w.synth.nz.mem[762] [5];
  assign _06948_ = \bapg_rd.w_ptr_r [1] ? _06947_ : _06946_;
  assign _06949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [5] : \MSYNC_1r1w.synth.nz.mem[764] [5];
  assign _06950_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [5] : \MSYNC_1r1w.synth.nz.mem[766] [5];
  assign _06951_ = \bapg_rd.w_ptr_r [1] ? _06950_ : _06949_;
  assign _06952_ = \bapg_rd.w_ptr_r [2] ? _06951_ : _06948_;
  assign _06953_ = \bapg_rd.w_ptr_r [3] ? _06952_ : _06945_;
  assign _06954_ = \bapg_rd.w_ptr_r [4] ? _06953_ : _06938_;
  assign _06955_ = \bapg_rd.w_ptr_r [5] ? _06954_ : _06923_;
  assign _06956_ = \bapg_rd.w_ptr_r [6] ? _06955_ : _06892_;
  assign _06957_ = \bapg_rd.w_ptr_r [7] ? _06956_ : _06829_;
  assign _06958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [5] : \MSYNC_1r1w.synth.nz.mem[768] [5];
  assign _06959_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [5] : \MSYNC_1r1w.synth.nz.mem[770] [5];
  assign _06960_ = \bapg_rd.w_ptr_r [1] ? _06959_ : _06958_;
  assign _06961_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [5] : \MSYNC_1r1w.synth.nz.mem[772] [5];
  assign _06962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [5] : \MSYNC_1r1w.synth.nz.mem[774] [5];
  assign _06963_ = \bapg_rd.w_ptr_r [1] ? _06962_ : _06961_;
  assign _06964_ = \bapg_rd.w_ptr_r [2] ? _06963_ : _06960_;
  assign _06965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [5] : \MSYNC_1r1w.synth.nz.mem[776] [5];
  assign _06966_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [5] : \MSYNC_1r1w.synth.nz.mem[778] [5];
  assign _06967_ = \bapg_rd.w_ptr_r [1] ? _06966_ : _06965_;
  assign _06968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [5] : \MSYNC_1r1w.synth.nz.mem[780] [5];
  assign _06969_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [5] : \MSYNC_1r1w.synth.nz.mem[782] [5];
  assign _06970_ = \bapg_rd.w_ptr_r [1] ? _06969_ : _06968_;
  assign _06971_ = \bapg_rd.w_ptr_r [2] ? _06970_ : _06967_;
  assign _06972_ = \bapg_rd.w_ptr_r [3] ? _06971_ : _06964_;
  assign _06973_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [5] : \MSYNC_1r1w.synth.nz.mem[784] [5];
  assign _06974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [5] : \MSYNC_1r1w.synth.nz.mem[786] [5];
  assign _06975_ = \bapg_rd.w_ptr_r [1] ? _06974_ : _06973_;
  assign _06976_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [5] : \MSYNC_1r1w.synth.nz.mem[788] [5];
  assign _06977_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [5] : \MSYNC_1r1w.synth.nz.mem[790] [5];
  assign _06978_ = \bapg_rd.w_ptr_r [1] ? _06977_ : _06976_;
  assign _06979_ = \bapg_rd.w_ptr_r [2] ? _06978_ : _06975_;
  assign _06980_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [5] : \MSYNC_1r1w.synth.nz.mem[792] [5];
  assign _06981_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [5] : \MSYNC_1r1w.synth.nz.mem[794] [5];
  assign _06982_ = \bapg_rd.w_ptr_r [1] ? _06981_ : _06980_;
  assign _06983_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [5] : \MSYNC_1r1w.synth.nz.mem[796] [5];
  assign _06984_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [5] : \MSYNC_1r1w.synth.nz.mem[798] [5];
  assign _06985_ = \bapg_rd.w_ptr_r [1] ? _06984_ : _06983_;
  assign _06986_ = \bapg_rd.w_ptr_r [2] ? _06985_ : _06982_;
  assign _06987_ = \bapg_rd.w_ptr_r [3] ? _06986_ : _06979_;
  assign _06988_ = \bapg_rd.w_ptr_r [4] ? _06987_ : _06972_;
  assign _06989_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [5] : \MSYNC_1r1w.synth.nz.mem[800] [5];
  assign _06990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [5] : \MSYNC_1r1w.synth.nz.mem[802] [5];
  assign _06991_ = \bapg_rd.w_ptr_r [1] ? _06990_ : _06989_;
  assign _06992_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [5] : \MSYNC_1r1w.synth.nz.mem[804] [5];
  assign _06993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [5] : \MSYNC_1r1w.synth.nz.mem[806] [5];
  assign _06994_ = \bapg_rd.w_ptr_r [1] ? _06993_ : _06992_;
  assign _06995_ = \bapg_rd.w_ptr_r [2] ? _06994_ : _06991_;
  assign _06996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [5] : \MSYNC_1r1w.synth.nz.mem[808] [5];
  assign _06997_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [5] : \MSYNC_1r1w.synth.nz.mem[810] [5];
  assign _06998_ = \bapg_rd.w_ptr_r [1] ? _06997_ : _06996_;
  assign _06999_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [5] : \MSYNC_1r1w.synth.nz.mem[812] [5];
  assign _07000_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [5] : \MSYNC_1r1w.synth.nz.mem[814] [5];
  assign _07001_ = \bapg_rd.w_ptr_r [1] ? _07000_ : _06999_;
  assign _07002_ = \bapg_rd.w_ptr_r [2] ? _07001_ : _06998_;
  assign _07003_ = \bapg_rd.w_ptr_r [3] ? _07002_ : _06995_;
  assign _07004_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [5] : \MSYNC_1r1w.synth.nz.mem[816] [5];
  assign _07005_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [5] : \MSYNC_1r1w.synth.nz.mem[818] [5];
  assign _07006_ = \bapg_rd.w_ptr_r [1] ? _07005_ : _07004_;
  assign _07007_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [5] : \MSYNC_1r1w.synth.nz.mem[820] [5];
  assign _07008_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [5] : \MSYNC_1r1w.synth.nz.mem[822] [5];
  assign _07009_ = \bapg_rd.w_ptr_r [1] ? _07008_ : _07007_;
  assign _07010_ = \bapg_rd.w_ptr_r [2] ? _07009_ : _07006_;
  assign _07011_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [5] : \MSYNC_1r1w.synth.nz.mem[824] [5];
  assign _07012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [5] : \MSYNC_1r1w.synth.nz.mem[826] [5];
  assign _07013_ = \bapg_rd.w_ptr_r [1] ? _07012_ : _07011_;
  assign _07014_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [5] : \MSYNC_1r1w.synth.nz.mem[828] [5];
  assign _07015_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [5] : \MSYNC_1r1w.synth.nz.mem[830] [5];
  assign _07016_ = \bapg_rd.w_ptr_r [1] ? _07015_ : _07014_;
  assign _07017_ = \bapg_rd.w_ptr_r [2] ? _07016_ : _07013_;
  assign _07018_ = \bapg_rd.w_ptr_r [3] ? _07017_ : _07010_;
  assign _07019_ = \bapg_rd.w_ptr_r [4] ? _07018_ : _07003_;
  assign _07020_ = \bapg_rd.w_ptr_r [5] ? _07019_ : _06988_;
  assign _07021_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [5] : \MSYNC_1r1w.synth.nz.mem[832] [5];
  assign _07022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [5] : \MSYNC_1r1w.synth.nz.mem[834] [5];
  assign _07023_ = \bapg_rd.w_ptr_r [1] ? _07022_ : _07021_;
  assign _07024_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [5] : \MSYNC_1r1w.synth.nz.mem[836] [5];
  assign _07025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [5] : \MSYNC_1r1w.synth.nz.mem[838] [5];
  assign _07026_ = \bapg_rd.w_ptr_r [1] ? _07025_ : _07024_;
  assign _07027_ = \bapg_rd.w_ptr_r [2] ? _07026_ : _07023_;
  assign _07028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [5] : \MSYNC_1r1w.synth.nz.mem[840] [5];
  assign _07029_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [5] : \MSYNC_1r1w.synth.nz.mem[842] [5];
  assign _07030_ = \bapg_rd.w_ptr_r [1] ? _07029_ : _07028_;
  assign _07031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [5] : \MSYNC_1r1w.synth.nz.mem[844] [5];
  assign _07032_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [5] : \MSYNC_1r1w.synth.nz.mem[846] [5];
  assign _07033_ = \bapg_rd.w_ptr_r [1] ? _07032_ : _07031_;
  assign _07034_ = \bapg_rd.w_ptr_r [2] ? _07033_ : _07030_;
  assign _07035_ = \bapg_rd.w_ptr_r [3] ? _07034_ : _07027_;
  assign _07036_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [5] : \MSYNC_1r1w.synth.nz.mem[848] [5];
  assign _07037_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [5] : \MSYNC_1r1w.synth.nz.mem[850] [5];
  assign _07038_ = \bapg_rd.w_ptr_r [1] ? _07037_ : _07036_;
  assign _07039_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [5] : \MSYNC_1r1w.synth.nz.mem[852] [5];
  assign _07040_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [5] : \MSYNC_1r1w.synth.nz.mem[854] [5];
  assign _07041_ = \bapg_rd.w_ptr_r [1] ? _07040_ : _07039_;
  assign _07042_ = \bapg_rd.w_ptr_r [2] ? _07041_ : _07038_;
  assign _07043_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [5] : \MSYNC_1r1w.synth.nz.mem[856] [5];
  assign _07044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [5] : \MSYNC_1r1w.synth.nz.mem[858] [5];
  assign _07045_ = \bapg_rd.w_ptr_r [1] ? _07044_ : _07043_;
  assign _07046_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [5] : \MSYNC_1r1w.synth.nz.mem[860] [5];
  assign _07047_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [5] : \MSYNC_1r1w.synth.nz.mem[862] [5];
  assign _07048_ = \bapg_rd.w_ptr_r [1] ? _07047_ : _07046_;
  assign _07049_ = \bapg_rd.w_ptr_r [2] ? _07048_ : _07045_;
  assign _07050_ = \bapg_rd.w_ptr_r [3] ? _07049_ : _07042_;
  assign _07051_ = \bapg_rd.w_ptr_r [4] ? _07050_ : _07035_;
  assign _07052_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [5] : \MSYNC_1r1w.synth.nz.mem[864] [5];
  assign _07053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [5] : \MSYNC_1r1w.synth.nz.mem[866] [5];
  assign _07054_ = \bapg_rd.w_ptr_r [1] ? _07053_ : _07052_;
  assign _07055_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [5] : \MSYNC_1r1w.synth.nz.mem[868] [5];
  assign _07056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [5] : \MSYNC_1r1w.synth.nz.mem[870] [5];
  assign _07057_ = \bapg_rd.w_ptr_r [1] ? _07056_ : _07055_;
  assign _07058_ = \bapg_rd.w_ptr_r [2] ? _07057_ : _07054_;
  assign _07059_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [5] : \MSYNC_1r1w.synth.nz.mem[872] [5];
  assign _07060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [5] : \MSYNC_1r1w.synth.nz.mem[874] [5];
  assign _07061_ = \bapg_rd.w_ptr_r [1] ? _07060_ : _07059_;
  assign _07062_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [5] : \MSYNC_1r1w.synth.nz.mem[876] [5];
  assign _07063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [5] : \MSYNC_1r1w.synth.nz.mem[878] [5];
  assign _07064_ = \bapg_rd.w_ptr_r [1] ? _07063_ : _07062_;
  assign _07065_ = \bapg_rd.w_ptr_r [2] ? _07064_ : _07061_;
  assign _07066_ = \bapg_rd.w_ptr_r [3] ? _07065_ : _07058_;
  assign _07067_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [5] : \MSYNC_1r1w.synth.nz.mem[880] [5];
  assign _07068_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [5] : \MSYNC_1r1w.synth.nz.mem[882] [5];
  assign _07069_ = \bapg_rd.w_ptr_r [1] ? _07068_ : _07067_;
  assign _07070_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [5] : \MSYNC_1r1w.synth.nz.mem[884] [5];
  assign _07071_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [5] : \MSYNC_1r1w.synth.nz.mem[886] [5];
  assign _07072_ = \bapg_rd.w_ptr_r [1] ? _07071_ : _07070_;
  assign _07073_ = \bapg_rd.w_ptr_r [2] ? _07072_ : _07069_;
  assign _07074_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [5] : \MSYNC_1r1w.synth.nz.mem[888] [5];
  assign _07075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [5] : \MSYNC_1r1w.synth.nz.mem[890] [5];
  assign _07076_ = \bapg_rd.w_ptr_r [1] ? _07075_ : _07074_;
  assign _07077_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [5] : \MSYNC_1r1w.synth.nz.mem[892] [5];
  assign _07078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [5] : \MSYNC_1r1w.synth.nz.mem[894] [5];
  assign _07079_ = \bapg_rd.w_ptr_r [1] ? _07078_ : _07077_;
  assign _07080_ = \bapg_rd.w_ptr_r [2] ? _07079_ : _07076_;
  assign _07081_ = \bapg_rd.w_ptr_r [3] ? _07080_ : _07073_;
  assign _07082_ = \bapg_rd.w_ptr_r [4] ? _07081_ : _07066_;
  assign _07083_ = \bapg_rd.w_ptr_r [5] ? _07082_ : _07051_;
  assign _07084_ = \bapg_rd.w_ptr_r [6] ? _07083_ : _07020_;
  assign _07085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [5] : \MSYNC_1r1w.synth.nz.mem[896] [5];
  assign _07086_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [5] : \MSYNC_1r1w.synth.nz.mem[898] [5];
  assign _07087_ = \bapg_rd.w_ptr_r [1] ? _07086_ : _07085_;
  assign _07088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [5] : \MSYNC_1r1w.synth.nz.mem[900] [5];
  assign _07089_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [5] : \MSYNC_1r1w.synth.nz.mem[902] [5];
  assign _07090_ = \bapg_rd.w_ptr_r [1] ? _07089_ : _07088_;
  assign _07091_ = \bapg_rd.w_ptr_r [2] ? _07090_ : _07087_;
  assign _07092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [5] : \MSYNC_1r1w.synth.nz.mem[904] [5];
  assign _07093_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [5] : \MSYNC_1r1w.synth.nz.mem[906] [5];
  assign _07094_ = \bapg_rd.w_ptr_r [1] ? _07093_ : _07092_;
  assign _07095_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [5] : \MSYNC_1r1w.synth.nz.mem[908] [5];
  assign _07096_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [5] : \MSYNC_1r1w.synth.nz.mem[910] [5];
  assign _07097_ = \bapg_rd.w_ptr_r [1] ? _07096_ : _07095_;
  assign _07098_ = \bapg_rd.w_ptr_r [2] ? _07097_ : _07094_;
  assign _07099_ = \bapg_rd.w_ptr_r [3] ? _07098_ : _07091_;
  assign _07100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [5] : \MSYNC_1r1w.synth.nz.mem[912] [5];
  assign _07101_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [5] : \MSYNC_1r1w.synth.nz.mem[914] [5];
  assign _07102_ = \bapg_rd.w_ptr_r [1] ? _07101_ : _07100_;
  assign _07103_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [5] : \MSYNC_1r1w.synth.nz.mem[916] [5];
  assign _07104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [5] : \MSYNC_1r1w.synth.nz.mem[918] [5];
  assign _07105_ = \bapg_rd.w_ptr_r [1] ? _07104_ : _07103_;
  assign _07106_ = \bapg_rd.w_ptr_r [2] ? _07105_ : _07102_;
  assign _07107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [5] : \MSYNC_1r1w.synth.nz.mem[920] [5];
  assign _07108_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [5] : \MSYNC_1r1w.synth.nz.mem[922] [5];
  assign _07109_ = \bapg_rd.w_ptr_r [1] ? _07108_ : _07107_;
  assign _07110_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [5] : \MSYNC_1r1w.synth.nz.mem[924] [5];
  assign _07111_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [5] : \MSYNC_1r1w.synth.nz.mem[926] [5];
  assign _07112_ = \bapg_rd.w_ptr_r [1] ? _07111_ : _07110_;
  assign _07113_ = \bapg_rd.w_ptr_r [2] ? _07112_ : _07109_;
  assign _07114_ = \bapg_rd.w_ptr_r [3] ? _07113_ : _07106_;
  assign _07115_ = \bapg_rd.w_ptr_r [4] ? _07114_ : _07099_;
  assign _07116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [5] : \MSYNC_1r1w.synth.nz.mem[928] [5];
  assign _07117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [5] : \MSYNC_1r1w.synth.nz.mem[930] [5];
  assign _07118_ = \bapg_rd.w_ptr_r [1] ? _07117_ : _07116_;
  assign _07119_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [5] : \MSYNC_1r1w.synth.nz.mem[932] [5];
  assign _07120_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [5] : \MSYNC_1r1w.synth.nz.mem[934] [5];
  assign _07121_ = \bapg_rd.w_ptr_r [1] ? _07120_ : _07119_;
  assign _07122_ = \bapg_rd.w_ptr_r [2] ? _07121_ : _07118_;
  assign _07123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [5] : \MSYNC_1r1w.synth.nz.mem[936] [5];
  assign _07124_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [5] : \MSYNC_1r1w.synth.nz.mem[938] [5];
  assign _07125_ = \bapg_rd.w_ptr_r [1] ? _07124_ : _07123_;
  assign _07126_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [5] : \MSYNC_1r1w.synth.nz.mem[940] [5];
  assign _07127_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [5] : \MSYNC_1r1w.synth.nz.mem[942] [5];
  assign _07128_ = \bapg_rd.w_ptr_r [1] ? _07127_ : _07126_;
  assign _07129_ = \bapg_rd.w_ptr_r [2] ? _07128_ : _07125_;
  assign _07130_ = \bapg_rd.w_ptr_r [3] ? _07129_ : _07122_;
  assign _07131_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [5] : \MSYNC_1r1w.synth.nz.mem[944] [5];
  assign _07132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [5] : \MSYNC_1r1w.synth.nz.mem[946] [5];
  assign _07133_ = \bapg_rd.w_ptr_r [1] ? _07132_ : _07131_;
  assign _07134_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [5] : \MSYNC_1r1w.synth.nz.mem[948] [5];
  assign _07135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [5] : \MSYNC_1r1w.synth.nz.mem[950] [5];
  assign _07136_ = \bapg_rd.w_ptr_r [1] ? _07135_ : _07134_;
  assign _07137_ = \bapg_rd.w_ptr_r [2] ? _07136_ : _07133_;
  assign _07138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [5] : \MSYNC_1r1w.synth.nz.mem[952] [5];
  assign _07139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [5] : \MSYNC_1r1w.synth.nz.mem[954] [5];
  assign _07140_ = \bapg_rd.w_ptr_r [1] ? _07139_ : _07138_;
  assign _07141_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [5] : \MSYNC_1r1w.synth.nz.mem[956] [5];
  assign _07142_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [5] : \MSYNC_1r1w.synth.nz.mem[958] [5];
  assign _07143_ = \bapg_rd.w_ptr_r [1] ? _07142_ : _07141_;
  assign _07144_ = \bapg_rd.w_ptr_r [2] ? _07143_ : _07140_;
  assign _07145_ = \bapg_rd.w_ptr_r [3] ? _07144_ : _07137_;
  assign _07146_ = \bapg_rd.w_ptr_r [4] ? _07145_ : _07130_;
  assign _07147_ = \bapg_rd.w_ptr_r [5] ? _07146_ : _07115_;
  assign _07148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [5] : \MSYNC_1r1w.synth.nz.mem[960] [5];
  assign _07149_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [5] : \MSYNC_1r1w.synth.nz.mem[962] [5];
  assign _07150_ = \bapg_rd.w_ptr_r [1] ? _07149_ : _07148_;
  assign _07151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [5] : \MSYNC_1r1w.synth.nz.mem[964] [5];
  assign _07152_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [5] : \MSYNC_1r1w.synth.nz.mem[966] [5];
  assign _07153_ = \bapg_rd.w_ptr_r [1] ? _07152_ : _07151_;
  assign _07154_ = \bapg_rd.w_ptr_r [2] ? _07153_ : _07150_;
  assign _07155_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [5] : \MSYNC_1r1w.synth.nz.mem[968] [5];
  assign _07156_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [5] : \MSYNC_1r1w.synth.nz.mem[970] [5];
  assign _07157_ = \bapg_rd.w_ptr_r [1] ? _07156_ : _07155_;
  assign _07158_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [5] : \MSYNC_1r1w.synth.nz.mem[972] [5];
  assign _07159_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [5] : \MSYNC_1r1w.synth.nz.mem[974] [5];
  assign _07160_ = \bapg_rd.w_ptr_r [1] ? _07159_ : _07158_;
  assign _07161_ = \bapg_rd.w_ptr_r [2] ? _07160_ : _07157_;
  assign _07162_ = \bapg_rd.w_ptr_r [3] ? _07161_ : _07154_;
  assign _07163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [5] : \MSYNC_1r1w.synth.nz.mem[976] [5];
  assign _07164_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [5] : \MSYNC_1r1w.synth.nz.mem[978] [5];
  assign _07165_ = \bapg_rd.w_ptr_r [1] ? _07164_ : _07163_;
  assign _07166_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [5] : \MSYNC_1r1w.synth.nz.mem[980] [5];
  assign _07167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [5] : \MSYNC_1r1w.synth.nz.mem[982] [5];
  assign _07168_ = \bapg_rd.w_ptr_r [1] ? _07167_ : _07166_;
  assign _07169_ = \bapg_rd.w_ptr_r [2] ? _07168_ : _07165_;
  assign _07170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [5] : \MSYNC_1r1w.synth.nz.mem[984] [5];
  assign _07171_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [5] : \MSYNC_1r1w.synth.nz.mem[986] [5];
  assign _07172_ = \bapg_rd.w_ptr_r [1] ? _07171_ : _07170_;
  assign _07173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [5] : \MSYNC_1r1w.synth.nz.mem[988] [5];
  assign _07174_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [5] : \MSYNC_1r1w.synth.nz.mem[990] [5];
  assign _07175_ = \bapg_rd.w_ptr_r [1] ? _07174_ : _07173_;
  assign _07176_ = \bapg_rd.w_ptr_r [2] ? _07175_ : _07172_;
  assign _07177_ = \bapg_rd.w_ptr_r [3] ? _07176_ : _07169_;
  assign _07178_ = \bapg_rd.w_ptr_r [4] ? _07177_ : _07162_;
  assign _07179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [5] : \MSYNC_1r1w.synth.nz.mem[992] [5];
  assign _07180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [5] : \MSYNC_1r1w.synth.nz.mem[994] [5];
  assign _07181_ = \bapg_rd.w_ptr_r [1] ? _07180_ : _07179_;
  assign _07182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [5] : \MSYNC_1r1w.synth.nz.mem[996] [5];
  assign _07183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [5] : \MSYNC_1r1w.synth.nz.mem[998] [5];
  assign _07184_ = \bapg_rd.w_ptr_r [1] ? _07183_ : _07182_;
  assign _07185_ = \bapg_rd.w_ptr_r [2] ? _07184_ : _07181_;
  assign _07186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [5] : \MSYNC_1r1w.synth.nz.mem[1000] [5];
  assign _07187_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [5] : \MSYNC_1r1w.synth.nz.mem[1002] [5];
  assign _07188_ = \bapg_rd.w_ptr_r [1] ? _07187_ : _07186_;
  assign _07189_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [5] : \MSYNC_1r1w.synth.nz.mem[1004] [5];
  assign _07190_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [5] : \MSYNC_1r1w.synth.nz.mem[1006] [5];
  assign _07191_ = \bapg_rd.w_ptr_r [1] ? _07190_ : _07189_;
  assign _07192_ = \bapg_rd.w_ptr_r [2] ? _07191_ : _07188_;
  assign _07193_ = \bapg_rd.w_ptr_r [3] ? _07192_ : _07185_;
  assign _07194_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [5] : \MSYNC_1r1w.synth.nz.mem[1008] [5];
  assign _07195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [5] : \MSYNC_1r1w.synth.nz.mem[1010] [5];
  assign _07196_ = \bapg_rd.w_ptr_r [1] ? _07195_ : _07194_;
  assign _07197_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [5] : \MSYNC_1r1w.synth.nz.mem[1012] [5];
  assign _07198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [5] : \MSYNC_1r1w.synth.nz.mem[1014] [5];
  assign _07199_ = \bapg_rd.w_ptr_r [1] ? _07198_ : _07197_;
  assign _07200_ = \bapg_rd.w_ptr_r [2] ? _07199_ : _07196_;
  assign _07201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [5] : \MSYNC_1r1w.synth.nz.mem[1016] [5];
  assign _07202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [5] : \MSYNC_1r1w.synth.nz.mem[1018] [5];
  assign _07203_ = \bapg_rd.w_ptr_r [1] ? _07202_ : _07201_;
  assign _07204_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [5] : \MSYNC_1r1w.synth.nz.mem[1020] [5];
  assign _07205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [5] : \MSYNC_1r1w.synth.nz.mem[1022] [5];
  assign _07206_ = \bapg_rd.w_ptr_r [1] ? _07205_ : _07204_;
  assign _07207_ = \bapg_rd.w_ptr_r [2] ? _07206_ : _07203_;
  assign _07208_ = \bapg_rd.w_ptr_r [3] ? _07207_ : _07200_;
  assign _07209_ = \bapg_rd.w_ptr_r [4] ? _07208_ : _07193_;
  assign _07210_ = \bapg_rd.w_ptr_r [5] ? _07209_ : _07178_;
  assign _07211_ = \bapg_rd.w_ptr_r [6] ? _07210_ : _07147_;
  assign _07212_ = \bapg_rd.w_ptr_r [7] ? _07211_ : _07084_;
  assign _07213_ = \bapg_rd.w_ptr_r [8] ? _07212_ : _06957_;
  assign r_data_o[5] = \bapg_rd.w_ptr_r [9] ? _07213_ : _06702_;
  assign _07214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [6] : \MSYNC_1r1w.synth.nz.mem[0] [6];
  assign _07215_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [6] : \MSYNC_1r1w.synth.nz.mem[2] [6];
  assign _07216_ = \bapg_rd.w_ptr_r [1] ? _07215_ : _07214_;
  assign _07217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [6] : \MSYNC_1r1w.synth.nz.mem[4] [6];
  assign _07218_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [6] : \MSYNC_1r1w.synth.nz.mem[6] [6];
  assign _07219_ = \bapg_rd.w_ptr_r [1] ? _07218_ : _07217_;
  assign _07220_ = \bapg_rd.w_ptr_r [2] ? _07219_ : _07216_;
  assign _07221_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [6] : \MSYNC_1r1w.synth.nz.mem[8] [6];
  assign _07222_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [6] : \MSYNC_1r1w.synth.nz.mem[10] [6];
  assign _07223_ = \bapg_rd.w_ptr_r [1] ? _07222_ : _07221_;
  assign _07224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [6] : \MSYNC_1r1w.synth.nz.mem[12] [6];
  assign _07225_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [6] : \MSYNC_1r1w.synth.nz.mem[14] [6];
  assign _07226_ = \bapg_rd.w_ptr_r [1] ? _07225_ : _07224_;
  assign _07227_ = \bapg_rd.w_ptr_r [2] ? _07226_ : _07223_;
  assign _07228_ = \bapg_rd.w_ptr_r [3] ? _07227_ : _07220_;
  assign _07229_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [6] : \MSYNC_1r1w.synth.nz.mem[16] [6];
  assign _07230_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [6] : \MSYNC_1r1w.synth.nz.mem[18] [6];
  assign _07231_ = \bapg_rd.w_ptr_r [1] ? _07230_ : _07229_;
  assign _07232_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [6] : \MSYNC_1r1w.synth.nz.mem[20] [6];
  assign _07233_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [6] : \MSYNC_1r1w.synth.nz.mem[22] [6];
  assign _07234_ = \bapg_rd.w_ptr_r [1] ? _07233_ : _07232_;
  assign _07235_ = \bapg_rd.w_ptr_r [2] ? _07234_ : _07231_;
  assign _07236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [6] : \MSYNC_1r1w.synth.nz.mem[24] [6];
  assign _07237_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [6] : \MSYNC_1r1w.synth.nz.mem[26] [6];
  assign _07238_ = \bapg_rd.w_ptr_r [1] ? _07237_ : _07236_;
  assign _07239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [6] : \MSYNC_1r1w.synth.nz.mem[28] [6];
  assign _07240_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [6] : \MSYNC_1r1w.synth.nz.mem[30] [6];
  assign _07241_ = \bapg_rd.w_ptr_r [1] ? _07240_ : _07239_;
  assign _07242_ = \bapg_rd.w_ptr_r [2] ? _07241_ : _07238_;
  assign _07243_ = \bapg_rd.w_ptr_r [3] ? _07242_ : _07235_;
  assign _07244_ = \bapg_rd.w_ptr_r [4] ? _07243_ : _07228_;
  assign _07245_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [6] : \MSYNC_1r1w.synth.nz.mem[32] [6];
  assign _07246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [6] : \MSYNC_1r1w.synth.nz.mem[34] [6];
  assign _07247_ = \bapg_rd.w_ptr_r [1] ? _07246_ : _07245_;
  assign _07248_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [6] : \MSYNC_1r1w.synth.nz.mem[36] [6];
  assign _07249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [6] : \MSYNC_1r1w.synth.nz.mem[38] [6];
  assign _07250_ = \bapg_rd.w_ptr_r [1] ? _07249_ : _07248_;
  assign _07251_ = \bapg_rd.w_ptr_r [2] ? _07250_ : _07247_;
  assign _07252_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [6] : \MSYNC_1r1w.synth.nz.mem[40] [6];
  assign _07253_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [6] : \MSYNC_1r1w.synth.nz.mem[42] [6];
  assign _07254_ = \bapg_rd.w_ptr_r [1] ? _07253_ : _07252_;
  assign _07255_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [6] : \MSYNC_1r1w.synth.nz.mem[44] [6];
  assign _07256_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [6] : \MSYNC_1r1w.synth.nz.mem[46] [6];
  assign _07257_ = \bapg_rd.w_ptr_r [1] ? _07256_ : _07255_;
  assign _07258_ = \bapg_rd.w_ptr_r [2] ? _07257_ : _07254_;
  assign _07259_ = \bapg_rd.w_ptr_r [3] ? _07258_ : _07251_;
  assign _07260_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [6] : \MSYNC_1r1w.synth.nz.mem[48] [6];
  assign _07261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [6] : \MSYNC_1r1w.synth.nz.mem[50] [6];
  assign _07262_ = \bapg_rd.w_ptr_r [1] ? _07261_ : _07260_;
  assign _07263_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [6] : \MSYNC_1r1w.synth.nz.mem[52] [6];
  assign _07264_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [6] : \MSYNC_1r1w.synth.nz.mem[54] [6];
  assign _07265_ = \bapg_rd.w_ptr_r [1] ? _07264_ : _07263_;
  assign _07266_ = \bapg_rd.w_ptr_r [2] ? _07265_ : _07262_;
  assign _07267_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [6] : \MSYNC_1r1w.synth.nz.mem[56] [6];
  assign _07268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [6] : \MSYNC_1r1w.synth.nz.mem[58] [6];
  assign _07269_ = \bapg_rd.w_ptr_r [1] ? _07268_ : _07267_;
  assign _07270_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [6] : \MSYNC_1r1w.synth.nz.mem[60] [6];
  assign _07271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [6] : \MSYNC_1r1w.synth.nz.mem[62] [6];
  assign _07272_ = \bapg_rd.w_ptr_r [1] ? _07271_ : _07270_;
  assign _07273_ = \bapg_rd.w_ptr_r [2] ? _07272_ : _07269_;
  assign _07274_ = \bapg_rd.w_ptr_r [3] ? _07273_ : _07266_;
  assign _07275_ = \bapg_rd.w_ptr_r [4] ? _07274_ : _07259_;
  assign _07276_ = \bapg_rd.w_ptr_r [5] ? _07275_ : _07244_;
  assign _07277_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [6] : \MSYNC_1r1w.synth.nz.mem[64] [6];
  assign _07278_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [6] : \MSYNC_1r1w.synth.nz.mem[66] [6];
  assign _07279_ = \bapg_rd.w_ptr_r [1] ? _07278_ : _07277_;
  assign _07280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [6] : \MSYNC_1r1w.synth.nz.mem[68] [6];
  assign _07281_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [6] : \MSYNC_1r1w.synth.nz.mem[70] [6];
  assign _07282_ = \bapg_rd.w_ptr_r [1] ? _07281_ : _07280_;
  assign _07283_ = \bapg_rd.w_ptr_r [2] ? _07282_ : _07279_;
  assign _07284_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [6] : \MSYNC_1r1w.synth.nz.mem[72] [6];
  assign _07285_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [6] : \MSYNC_1r1w.synth.nz.mem[74] [6];
  assign _07286_ = \bapg_rd.w_ptr_r [1] ? _07285_ : _07284_;
  assign _07287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [6] : \MSYNC_1r1w.synth.nz.mem[76] [6];
  assign _07288_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [6] : \MSYNC_1r1w.synth.nz.mem[78] [6];
  assign _07289_ = \bapg_rd.w_ptr_r [1] ? _07288_ : _07287_;
  assign _07290_ = \bapg_rd.w_ptr_r [2] ? _07289_ : _07286_;
  assign _07291_ = \bapg_rd.w_ptr_r [3] ? _07290_ : _07283_;
  assign _07292_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [6] : \MSYNC_1r1w.synth.nz.mem[80] [6];
  assign _07293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [6] : \MSYNC_1r1w.synth.nz.mem[82] [6];
  assign _07294_ = \bapg_rd.w_ptr_r [1] ? _07293_ : _07292_;
  assign _07295_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [6] : \MSYNC_1r1w.synth.nz.mem[84] [6];
  assign _07296_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [6] : \MSYNC_1r1w.synth.nz.mem[86] [6];
  assign _07297_ = \bapg_rd.w_ptr_r [1] ? _07296_ : _07295_;
  assign _07298_ = \bapg_rd.w_ptr_r [2] ? _07297_ : _07294_;
  assign _07299_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [6] : \MSYNC_1r1w.synth.nz.mem[88] [6];
  assign _07300_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [6] : \MSYNC_1r1w.synth.nz.mem[90] [6];
  assign _07301_ = \bapg_rd.w_ptr_r [1] ? _07300_ : _07299_;
  assign _07302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [6] : \MSYNC_1r1w.synth.nz.mem[92] [6];
  assign _07303_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [6] : \MSYNC_1r1w.synth.nz.mem[94] [6];
  assign _07304_ = \bapg_rd.w_ptr_r [1] ? _07303_ : _07302_;
  assign _07305_ = \bapg_rd.w_ptr_r [2] ? _07304_ : _07301_;
  assign _07306_ = \bapg_rd.w_ptr_r [3] ? _07305_ : _07298_;
  assign _07307_ = \bapg_rd.w_ptr_r [4] ? _07306_ : _07291_;
  assign _07308_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [6] : \MSYNC_1r1w.synth.nz.mem[96] [6];
  assign _07309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [6] : \MSYNC_1r1w.synth.nz.mem[98] [6];
  assign _07310_ = \bapg_rd.w_ptr_r [1] ? _07309_ : _07308_;
  assign _07311_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [6] : \MSYNC_1r1w.synth.nz.mem[100] [6];
  assign _07312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [6] : \MSYNC_1r1w.synth.nz.mem[102] [6];
  assign _07313_ = \bapg_rd.w_ptr_r [1] ? _07312_ : _07311_;
  assign _07314_ = \bapg_rd.w_ptr_r [2] ? _07313_ : _07310_;
  assign _07315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [6] : \MSYNC_1r1w.synth.nz.mem[104] [6];
  assign _07316_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [6] : \MSYNC_1r1w.synth.nz.mem[106] [6];
  assign _07317_ = \bapg_rd.w_ptr_r [1] ? _07316_ : _07315_;
  assign _07318_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [6] : \MSYNC_1r1w.synth.nz.mem[108] [6];
  assign _07319_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [6] : \MSYNC_1r1w.synth.nz.mem[110] [6];
  assign _07320_ = \bapg_rd.w_ptr_r [1] ? _07319_ : _07318_;
  assign _07321_ = \bapg_rd.w_ptr_r [2] ? _07320_ : _07317_;
  assign _07322_ = \bapg_rd.w_ptr_r [3] ? _07321_ : _07314_;
  assign _07323_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [6] : \MSYNC_1r1w.synth.nz.mem[112] [6];
  assign _07324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [6] : \MSYNC_1r1w.synth.nz.mem[114] [6];
  assign _07325_ = \bapg_rd.w_ptr_r [1] ? _07324_ : _07323_;
  assign _07326_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [6] : \MSYNC_1r1w.synth.nz.mem[116] [6];
  assign _07327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [6] : \MSYNC_1r1w.synth.nz.mem[118] [6];
  assign _07328_ = \bapg_rd.w_ptr_r [1] ? _07327_ : _07326_;
  assign _07329_ = \bapg_rd.w_ptr_r [2] ? _07328_ : _07325_;
  assign _07330_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [6] : \MSYNC_1r1w.synth.nz.mem[120] [6];
  assign _07331_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [6] : \MSYNC_1r1w.synth.nz.mem[122] [6];
  assign _07332_ = \bapg_rd.w_ptr_r [1] ? _07331_ : _07330_;
  assign _07333_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [6] : \MSYNC_1r1w.synth.nz.mem[124] [6];
  assign _07334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [6] : \MSYNC_1r1w.synth.nz.mem[126] [6];
  assign _07335_ = \bapg_rd.w_ptr_r [1] ? _07334_ : _07333_;
  assign _07336_ = \bapg_rd.w_ptr_r [2] ? _07335_ : _07332_;
  assign _07337_ = \bapg_rd.w_ptr_r [3] ? _07336_ : _07329_;
  assign _07338_ = \bapg_rd.w_ptr_r [4] ? _07337_ : _07322_;
  assign _07339_ = \bapg_rd.w_ptr_r [5] ? _07338_ : _07307_;
  assign _07340_ = \bapg_rd.w_ptr_r [6] ? _07339_ : _07276_;
  assign _07341_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [6] : \MSYNC_1r1w.synth.nz.mem[128] [6];
  assign _07342_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [6] : \MSYNC_1r1w.synth.nz.mem[130] [6];
  assign _07343_ = \bapg_rd.w_ptr_r [1] ? _07342_ : _07341_;
  assign _07344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [6] : \MSYNC_1r1w.synth.nz.mem[132] [6];
  assign _07345_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [6] : \MSYNC_1r1w.synth.nz.mem[134] [6];
  assign _07346_ = \bapg_rd.w_ptr_r [1] ? _07345_ : _07344_;
  assign _07347_ = \bapg_rd.w_ptr_r [2] ? _07346_ : _07343_;
  assign _07348_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [6] : \MSYNC_1r1w.synth.nz.mem[136] [6];
  assign _07349_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [6] : \MSYNC_1r1w.synth.nz.mem[138] [6];
  assign _07350_ = \bapg_rd.w_ptr_r [1] ? _07349_ : _07348_;
  assign _07351_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [6] : \MSYNC_1r1w.synth.nz.mem[140] [6];
  assign _07352_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [6] : \MSYNC_1r1w.synth.nz.mem[142] [6];
  assign _07353_ = \bapg_rd.w_ptr_r [1] ? _07352_ : _07351_;
  assign _07354_ = \bapg_rd.w_ptr_r [2] ? _07353_ : _07350_;
  assign _07355_ = \bapg_rd.w_ptr_r [3] ? _07354_ : _07347_;
  assign _07356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [6] : \MSYNC_1r1w.synth.nz.mem[144] [6];
  assign _07357_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [6] : \MSYNC_1r1w.synth.nz.mem[146] [6];
  assign _07358_ = \bapg_rd.w_ptr_r [1] ? _07357_ : _07356_;
  assign _07359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [6] : \MSYNC_1r1w.synth.nz.mem[148] [6];
  assign _07360_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [6] : \MSYNC_1r1w.synth.nz.mem[150] [6];
  assign _07361_ = \bapg_rd.w_ptr_r [1] ? _07360_ : _07359_;
  assign _07362_ = \bapg_rd.w_ptr_r [2] ? _07361_ : _07358_;
  assign _07363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [6] : \MSYNC_1r1w.synth.nz.mem[152] [6];
  assign _07364_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [6] : \MSYNC_1r1w.synth.nz.mem[154] [6];
  assign _07365_ = \bapg_rd.w_ptr_r [1] ? _07364_ : _07363_;
  assign _07366_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [6] : \MSYNC_1r1w.synth.nz.mem[156] [6];
  assign _07367_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [6] : \MSYNC_1r1w.synth.nz.mem[158] [6];
  assign _07368_ = \bapg_rd.w_ptr_r [1] ? _07367_ : _07366_;
  assign _07369_ = \bapg_rd.w_ptr_r [2] ? _07368_ : _07365_;
  assign _07370_ = \bapg_rd.w_ptr_r [3] ? _07369_ : _07362_;
  assign _07371_ = \bapg_rd.w_ptr_r [4] ? _07370_ : _07355_;
  assign _07372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [6] : \MSYNC_1r1w.synth.nz.mem[160] [6];
  assign _07373_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [6] : \MSYNC_1r1w.synth.nz.mem[162] [6];
  assign _07374_ = \bapg_rd.w_ptr_r [1] ? _07373_ : _07372_;
  assign _07375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [6] : \MSYNC_1r1w.synth.nz.mem[164] [6];
  assign _07376_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [6] : \MSYNC_1r1w.synth.nz.mem[166] [6];
  assign _07377_ = \bapg_rd.w_ptr_r [1] ? _07376_ : _07375_;
  assign _07378_ = \bapg_rd.w_ptr_r [2] ? _07377_ : _07374_;
  assign _07379_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [6] : \MSYNC_1r1w.synth.nz.mem[168] [6];
  assign _07380_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [6] : \MSYNC_1r1w.synth.nz.mem[170] [6];
  assign _07381_ = \bapg_rd.w_ptr_r [1] ? _07380_ : _07379_;
  assign _07382_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [6] : \MSYNC_1r1w.synth.nz.mem[172] [6];
  assign _07383_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [6] : \MSYNC_1r1w.synth.nz.mem[174] [6];
  assign _07384_ = \bapg_rd.w_ptr_r [1] ? _07383_ : _07382_;
  assign _07385_ = \bapg_rd.w_ptr_r [2] ? _07384_ : _07381_;
  assign _07386_ = \bapg_rd.w_ptr_r [3] ? _07385_ : _07378_;
  assign _07387_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [6] : \MSYNC_1r1w.synth.nz.mem[176] [6];
  assign _07388_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [6] : \MSYNC_1r1w.synth.nz.mem[178] [6];
  assign _07389_ = \bapg_rd.w_ptr_r [1] ? _07388_ : _07387_;
  assign _07390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [6] : \MSYNC_1r1w.synth.nz.mem[180] [6];
  assign _07391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [6] : \MSYNC_1r1w.synth.nz.mem[182] [6];
  assign _07392_ = \bapg_rd.w_ptr_r [1] ? _07391_ : _07390_;
  assign _07393_ = \bapg_rd.w_ptr_r [2] ? _07392_ : _07389_;
  assign _07394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [6] : \MSYNC_1r1w.synth.nz.mem[184] [6];
  assign _07395_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [6] : \MSYNC_1r1w.synth.nz.mem[186] [6];
  assign _07396_ = \bapg_rd.w_ptr_r [1] ? _07395_ : _07394_;
  assign _07397_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [6] : \MSYNC_1r1w.synth.nz.mem[188] [6];
  assign _07398_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [6] : \MSYNC_1r1w.synth.nz.mem[190] [6];
  assign _07399_ = \bapg_rd.w_ptr_r [1] ? _07398_ : _07397_;
  assign _07400_ = \bapg_rd.w_ptr_r [2] ? _07399_ : _07396_;
  assign _07401_ = \bapg_rd.w_ptr_r [3] ? _07400_ : _07393_;
  assign _07402_ = \bapg_rd.w_ptr_r [4] ? _07401_ : _07386_;
  assign _07403_ = \bapg_rd.w_ptr_r [5] ? _07402_ : _07371_;
  assign _07404_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [6] : \MSYNC_1r1w.synth.nz.mem[192] [6];
  assign _07405_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [6] : \MSYNC_1r1w.synth.nz.mem[194] [6];
  assign _07406_ = \bapg_rd.w_ptr_r [1] ? _07405_ : _07404_;
  assign _07407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [6] : \MSYNC_1r1w.synth.nz.mem[196] [6];
  assign _07408_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [6] : \MSYNC_1r1w.synth.nz.mem[198] [6];
  assign _07409_ = \bapg_rd.w_ptr_r [1] ? _07408_ : _07407_;
  assign _07410_ = \bapg_rd.w_ptr_r [2] ? _07409_ : _07406_;
  assign _07411_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [6] : \MSYNC_1r1w.synth.nz.mem[200] [6];
  assign _07412_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [6] : \MSYNC_1r1w.synth.nz.mem[202] [6];
  assign _07413_ = \bapg_rd.w_ptr_r [1] ? _07412_ : _07411_;
  assign _07414_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [6] : \MSYNC_1r1w.synth.nz.mem[204] [6];
  assign _07415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [6] : \MSYNC_1r1w.synth.nz.mem[206] [6];
  assign _07416_ = \bapg_rd.w_ptr_r [1] ? _07415_ : _07414_;
  assign _07417_ = \bapg_rd.w_ptr_r [2] ? _07416_ : _07413_;
  assign _07418_ = \bapg_rd.w_ptr_r [3] ? _07417_ : _07410_;
  assign _07419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [6] : \MSYNC_1r1w.synth.nz.mem[208] [6];
  assign _07420_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [6] : \MSYNC_1r1w.synth.nz.mem[210] [6];
  assign _07421_ = \bapg_rd.w_ptr_r [1] ? _07420_ : _07419_;
  assign _07422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [6] : \MSYNC_1r1w.synth.nz.mem[212] [6];
  assign _07423_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [6] : \MSYNC_1r1w.synth.nz.mem[214] [6];
  assign _07424_ = \bapg_rd.w_ptr_r [1] ? _07423_ : _07422_;
  assign _07425_ = \bapg_rd.w_ptr_r [2] ? _07424_ : _07421_;
  assign _07426_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [6] : \MSYNC_1r1w.synth.nz.mem[216] [6];
  assign _07427_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [6] : \MSYNC_1r1w.synth.nz.mem[218] [6];
  assign _07428_ = \bapg_rd.w_ptr_r [1] ? _07427_ : _07426_;
  assign _07429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [6] : \MSYNC_1r1w.synth.nz.mem[220] [6];
  assign _07430_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [6] : \MSYNC_1r1w.synth.nz.mem[222] [6];
  assign _07431_ = \bapg_rd.w_ptr_r [1] ? _07430_ : _07429_;
  assign _07432_ = \bapg_rd.w_ptr_r [2] ? _07431_ : _07428_;
  assign _07433_ = \bapg_rd.w_ptr_r [3] ? _07432_ : _07425_;
  assign _07434_ = \bapg_rd.w_ptr_r [4] ? _07433_ : _07418_;
  assign _07435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [6] : \MSYNC_1r1w.synth.nz.mem[224] [6];
  assign _07436_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [6] : \MSYNC_1r1w.synth.nz.mem[226] [6];
  assign _07437_ = \bapg_rd.w_ptr_r [1] ? _07436_ : _07435_;
  assign _07438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [6] : \MSYNC_1r1w.synth.nz.mem[228] [6];
  assign _07439_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [6] : \MSYNC_1r1w.synth.nz.mem[230] [6];
  assign _07440_ = \bapg_rd.w_ptr_r [1] ? _07439_ : _07438_;
  assign _07441_ = \bapg_rd.w_ptr_r [2] ? _07440_ : _07437_;
  assign _07442_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [6] : \MSYNC_1r1w.synth.nz.mem[232] [6];
  assign _07443_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [6] : \MSYNC_1r1w.synth.nz.mem[234] [6];
  assign _07444_ = \bapg_rd.w_ptr_r [1] ? _07443_ : _07442_;
  assign _07445_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [6] : \MSYNC_1r1w.synth.nz.mem[236] [6];
  assign _07446_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [6] : \MSYNC_1r1w.synth.nz.mem[238] [6];
  assign _07447_ = \bapg_rd.w_ptr_r [1] ? _07446_ : _07445_;
  assign _07448_ = \bapg_rd.w_ptr_r [2] ? _07447_ : _07444_;
  assign _07449_ = \bapg_rd.w_ptr_r [3] ? _07448_ : _07441_;
  assign _07450_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [6] : \MSYNC_1r1w.synth.nz.mem[240] [6];
  assign _07451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [6] : \MSYNC_1r1w.synth.nz.mem[242] [6];
  assign _07452_ = \bapg_rd.w_ptr_r [1] ? _07451_ : _07450_;
  assign _07453_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [6] : \MSYNC_1r1w.synth.nz.mem[244] [6];
  assign _07454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [6] : \MSYNC_1r1w.synth.nz.mem[246] [6];
  assign _07455_ = \bapg_rd.w_ptr_r [1] ? _07454_ : _07453_;
  assign _07456_ = \bapg_rd.w_ptr_r [2] ? _07455_ : _07452_;
  assign _07457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [6] : \MSYNC_1r1w.synth.nz.mem[248] [6];
  assign _07458_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [6] : \MSYNC_1r1w.synth.nz.mem[250] [6];
  assign _07459_ = \bapg_rd.w_ptr_r [1] ? _07458_ : _07457_;
  assign _07460_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [6] : \MSYNC_1r1w.synth.nz.mem[252] [6];
  assign _07461_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [6] : \MSYNC_1r1w.synth.nz.mem[254] [6];
  assign _07462_ = \bapg_rd.w_ptr_r [1] ? _07461_ : _07460_;
  assign _07463_ = \bapg_rd.w_ptr_r [2] ? _07462_ : _07459_;
  assign _07464_ = \bapg_rd.w_ptr_r [3] ? _07463_ : _07456_;
  assign _07465_ = \bapg_rd.w_ptr_r [4] ? _07464_ : _07449_;
  assign _07466_ = \bapg_rd.w_ptr_r [5] ? _07465_ : _07434_;
  assign _07467_ = \bapg_rd.w_ptr_r [6] ? _07466_ : _07403_;
  assign _07468_ = \bapg_rd.w_ptr_r [7] ? _07467_ : _07340_;
  assign _07469_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [6] : \MSYNC_1r1w.synth.nz.mem[256] [6];
  assign _07470_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [6] : \MSYNC_1r1w.synth.nz.mem[258] [6];
  assign _07471_ = \bapg_rd.w_ptr_r [1] ? _07470_ : _07469_;
  assign _07472_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [6] : \MSYNC_1r1w.synth.nz.mem[260] [6];
  assign _07473_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [6] : \MSYNC_1r1w.synth.nz.mem[262] [6];
  assign _07474_ = \bapg_rd.w_ptr_r [1] ? _07473_ : _07472_;
  assign _07475_ = \bapg_rd.w_ptr_r [2] ? _07474_ : _07471_;
  assign _07476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [6] : \MSYNC_1r1w.synth.nz.mem[264] [6];
  assign _07477_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [6] : \MSYNC_1r1w.synth.nz.mem[266] [6];
  assign _07478_ = \bapg_rd.w_ptr_r [1] ? _07477_ : _07476_;
  assign _07479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [6] : \MSYNC_1r1w.synth.nz.mem[268] [6];
  assign _07480_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [6] : \MSYNC_1r1w.synth.nz.mem[270] [6];
  assign _07481_ = \bapg_rd.w_ptr_r [1] ? _07480_ : _07479_;
  assign _07482_ = \bapg_rd.w_ptr_r [2] ? _07481_ : _07478_;
  assign _07483_ = \bapg_rd.w_ptr_r [3] ? _07482_ : _07475_;
  assign _07484_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [6] : \MSYNC_1r1w.synth.nz.mem[272] [6];
  assign _07485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [6] : \MSYNC_1r1w.synth.nz.mem[274] [6];
  assign _07486_ = \bapg_rd.w_ptr_r [1] ? _07485_ : _07484_;
  assign _07487_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [6] : \MSYNC_1r1w.synth.nz.mem[276] [6];
  assign _07488_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [6] : \MSYNC_1r1w.synth.nz.mem[278] [6];
  assign _07489_ = \bapg_rd.w_ptr_r [1] ? _07488_ : _07487_;
  assign _07490_ = \bapg_rd.w_ptr_r [2] ? _07489_ : _07486_;
  assign _07491_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [6] : \MSYNC_1r1w.synth.nz.mem[280] [6];
  assign _07492_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [6] : \MSYNC_1r1w.synth.nz.mem[282] [6];
  assign _07493_ = \bapg_rd.w_ptr_r [1] ? _07492_ : _07491_;
  assign _07494_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [6] : \MSYNC_1r1w.synth.nz.mem[284] [6];
  assign _07495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [6] : \MSYNC_1r1w.synth.nz.mem[286] [6];
  assign _07496_ = \bapg_rd.w_ptr_r [1] ? _07495_ : _07494_;
  assign _07497_ = \bapg_rd.w_ptr_r [2] ? _07496_ : _07493_;
  assign _07498_ = \bapg_rd.w_ptr_r [3] ? _07497_ : _07490_;
  assign _07499_ = \bapg_rd.w_ptr_r [4] ? _07498_ : _07483_;
  assign _07500_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [6] : \MSYNC_1r1w.synth.nz.mem[288] [6];
  assign _07501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [6] : \MSYNC_1r1w.synth.nz.mem[290] [6];
  assign _07502_ = \bapg_rd.w_ptr_r [1] ? _07501_ : _07500_;
  assign _07503_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [6] : \MSYNC_1r1w.synth.nz.mem[292] [6];
  assign _07504_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [6] : \MSYNC_1r1w.synth.nz.mem[294] [6];
  assign _07505_ = \bapg_rd.w_ptr_r [1] ? _07504_ : _07503_;
  assign _07506_ = \bapg_rd.w_ptr_r [2] ? _07505_ : _07502_;
  assign _07507_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [6] : \MSYNC_1r1w.synth.nz.mem[296] [6];
  assign _07508_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [6] : \MSYNC_1r1w.synth.nz.mem[298] [6];
  assign _07509_ = \bapg_rd.w_ptr_r [1] ? _07508_ : _07507_;
  assign _07510_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [6] : \MSYNC_1r1w.synth.nz.mem[300] [6];
  assign _07511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [6] : \MSYNC_1r1w.synth.nz.mem[302] [6];
  assign _07512_ = \bapg_rd.w_ptr_r [1] ? _07511_ : _07510_;
  assign _07513_ = \bapg_rd.w_ptr_r [2] ? _07512_ : _07509_;
  assign _07514_ = \bapg_rd.w_ptr_r [3] ? _07513_ : _07506_;
  assign _07515_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [6] : \MSYNC_1r1w.synth.nz.mem[304] [6];
  assign _07516_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [6] : \MSYNC_1r1w.synth.nz.mem[306] [6];
  assign _07517_ = \bapg_rd.w_ptr_r [1] ? _07516_ : _07515_;
  assign _07518_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [6] : \MSYNC_1r1w.synth.nz.mem[308] [6];
  assign _07519_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [6] : \MSYNC_1r1w.synth.nz.mem[310] [6];
  assign _07520_ = \bapg_rd.w_ptr_r [1] ? _07519_ : _07518_;
  assign _07521_ = \bapg_rd.w_ptr_r [2] ? _07520_ : _07517_;
  assign _07522_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [6] : \MSYNC_1r1w.synth.nz.mem[312] [6];
  assign _07523_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [6] : \MSYNC_1r1w.synth.nz.mem[314] [6];
  assign _07524_ = \bapg_rd.w_ptr_r [1] ? _07523_ : _07522_;
  assign _07525_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [6] : \MSYNC_1r1w.synth.nz.mem[316] [6];
  assign _07526_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [6] : \MSYNC_1r1w.synth.nz.mem[318] [6];
  assign _07527_ = \bapg_rd.w_ptr_r [1] ? _07526_ : _07525_;
  assign _07528_ = \bapg_rd.w_ptr_r [2] ? _07527_ : _07524_;
  assign _07529_ = \bapg_rd.w_ptr_r [3] ? _07528_ : _07521_;
  assign _07530_ = \bapg_rd.w_ptr_r [4] ? _07529_ : _07514_;
  assign _07531_ = \bapg_rd.w_ptr_r [5] ? _07530_ : _07499_;
  assign _07532_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [6] : \MSYNC_1r1w.synth.nz.mem[320] [6];
  assign _07533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [6] : \MSYNC_1r1w.synth.nz.mem[322] [6];
  assign _07534_ = \bapg_rd.w_ptr_r [1] ? _07533_ : _07532_;
  assign _07535_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [6] : \MSYNC_1r1w.synth.nz.mem[324] [6];
  assign _07536_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [6] : \MSYNC_1r1w.synth.nz.mem[326] [6];
  assign _07537_ = \bapg_rd.w_ptr_r [1] ? _07536_ : _07535_;
  assign _07538_ = \bapg_rd.w_ptr_r [2] ? _07537_ : _07534_;
  assign _07539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [6] : \MSYNC_1r1w.synth.nz.mem[328] [6];
  assign _07540_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [6] : \MSYNC_1r1w.synth.nz.mem[330] [6];
  assign _07541_ = \bapg_rd.w_ptr_r [1] ? _07540_ : _07539_;
  assign _07542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [6] : \MSYNC_1r1w.synth.nz.mem[332] [6];
  assign _07543_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [6] : \MSYNC_1r1w.synth.nz.mem[334] [6];
  assign _07544_ = \bapg_rd.w_ptr_r [1] ? _07543_ : _07542_;
  assign _07545_ = \bapg_rd.w_ptr_r [2] ? _07544_ : _07541_;
  assign _07546_ = \bapg_rd.w_ptr_r [3] ? _07545_ : _07538_;
  assign _07547_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [6] : \MSYNC_1r1w.synth.nz.mem[336] [6];
  assign _07548_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [6] : \MSYNC_1r1w.synth.nz.mem[338] [6];
  assign _07549_ = \bapg_rd.w_ptr_r [1] ? _07548_ : _07547_;
  assign _07550_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [6] : \MSYNC_1r1w.synth.nz.mem[340] [6];
  assign _07551_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [6] : \MSYNC_1r1w.synth.nz.mem[342] [6];
  assign _07552_ = \bapg_rd.w_ptr_r [1] ? _07551_ : _07550_;
  assign _07553_ = \bapg_rd.w_ptr_r [2] ? _07552_ : _07549_;
  assign _07554_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [6] : \MSYNC_1r1w.synth.nz.mem[344] [6];
  assign _07555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [6] : \MSYNC_1r1w.synth.nz.mem[346] [6];
  assign _07556_ = \bapg_rd.w_ptr_r [1] ? _07555_ : _07554_;
  assign _07557_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [6] : \MSYNC_1r1w.synth.nz.mem[348] [6];
  assign _07558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [6] : \MSYNC_1r1w.synth.nz.mem[350] [6];
  assign _07559_ = \bapg_rd.w_ptr_r [1] ? _07558_ : _07557_;
  assign _07560_ = \bapg_rd.w_ptr_r [2] ? _07559_ : _07556_;
  assign _07561_ = \bapg_rd.w_ptr_r [3] ? _07560_ : _07553_;
  assign _07562_ = \bapg_rd.w_ptr_r [4] ? _07561_ : _07546_;
  assign _07563_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [6] : \MSYNC_1r1w.synth.nz.mem[352] [6];
  assign _07564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [6] : \MSYNC_1r1w.synth.nz.mem[354] [6];
  assign _07565_ = \bapg_rd.w_ptr_r [1] ? _07564_ : _07563_;
  assign _07566_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [6] : \MSYNC_1r1w.synth.nz.mem[356] [6];
  assign _07567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [6] : \MSYNC_1r1w.synth.nz.mem[358] [6];
  assign _07568_ = \bapg_rd.w_ptr_r [1] ? _07567_ : _07566_;
  assign _07569_ = \bapg_rd.w_ptr_r [2] ? _07568_ : _07565_;
  assign _07570_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [6] : \MSYNC_1r1w.synth.nz.mem[360] [6];
  assign _07571_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [6] : \MSYNC_1r1w.synth.nz.mem[362] [6];
  assign _07572_ = \bapg_rd.w_ptr_r [1] ? _07571_ : _07570_;
  assign _07573_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [6] : \MSYNC_1r1w.synth.nz.mem[364] [6];
  assign _07574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [6] : \MSYNC_1r1w.synth.nz.mem[366] [6];
  assign _07575_ = \bapg_rd.w_ptr_r [1] ? _07574_ : _07573_;
  assign _07576_ = \bapg_rd.w_ptr_r [2] ? _07575_ : _07572_;
  assign _07577_ = \bapg_rd.w_ptr_r [3] ? _07576_ : _07569_;
  assign _07578_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [6] : \MSYNC_1r1w.synth.nz.mem[368] [6];
  assign _07579_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [6] : \MSYNC_1r1w.synth.nz.mem[370] [6];
  assign _07580_ = \bapg_rd.w_ptr_r [1] ? _07579_ : _07578_;
  assign _07581_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [6] : \MSYNC_1r1w.synth.nz.mem[372] [6];
  assign _07582_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [6] : \MSYNC_1r1w.synth.nz.mem[374] [6];
  assign _07583_ = \bapg_rd.w_ptr_r [1] ? _07582_ : _07581_;
  assign _07584_ = \bapg_rd.w_ptr_r [2] ? _07583_ : _07580_;
  assign _07585_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [6] : \MSYNC_1r1w.synth.nz.mem[376] [6];
  assign _07586_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [6] : \MSYNC_1r1w.synth.nz.mem[378] [6];
  assign _07587_ = \bapg_rd.w_ptr_r [1] ? _07586_ : _07585_;
  assign _07588_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [6] : \MSYNC_1r1w.synth.nz.mem[380] [6];
  assign _07589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [6] : \MSYNC_1r1w.synth.nz.mem[382] [6];
  assign _07590_ = \bapg_rd.w_ptr_r [1] ? _07589_ : _07588_;
  assign _07591_ = \bapg_rd.w_ptr_r [2] ? _07590_ : _07587_;
  assign _07592_ = \bapg_rd.w_ptr_r [3] ? _07591_ : _07584_;
  assign _07593_ = \bapg_rd.w_ptr_r [4] ? _07592_ : _07577_;
  assign _07594_ = \bapg_rd.w_ptr_r [5] ? _07593_ : _07562_;
  assign _07595_ = \bapg_rd.w_ptr_r [6] ? _07594_ : _07531_;
  assign _07596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [6] : \MSYNC_1r1w.synth.nz.mem[384] [6];
  assign _07597_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [6] : \MSYNC_1r1w.synth.nz.mem[386] [6];
  assign _07598_ = \bapg_rd.w_ptr_r [1] ? _07597_ : _07596_;
  assign _07599_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [6] : \MSYNC_1r1w.synth.nz.mem[388] [6];
  assign _07600_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [6] : \MSYNC_1r1w.synth.nz.mem[390] [6];
  assign _07601_ = \bapg_rd.w_ptr_r [1] ? _07600_ : _07599_;
  assign _07602_ = \bapg_rd.w_ptr_r [2] ? _07601_ : _07598_;
  assign _07603_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [6] : \MSYNC_1r1w.synth.nz.mem[392] [6];
  assign _07604_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [6] : \MSYNC_1r1w.synth.nz.mem[394] [6];
  assign _07605_ = \bapg_rd.w_ptr_r [1] ? _07604_ : _07603_;
  assign _07606_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [6] : \MSYNC_1r1w.synth.nz.mem[396] [6];
  assign _07607_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [6] : \MSYNC_1r1w.synth.nz.mem[398] [6];
  assign _07608_ = \bapg_rd.w_ptr_r [1] ? _07607_ : _07606_;
  assign _07609_ = \bapg_rd.w_ptr_r [2] ? _07608_ : _07605_;
  assign _07610_ = \bapg_rd.w_ptr_r [3] ? _07609_ : _07602_;
  assign _07611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [6] : \MSYNC_1r1w.synth.nz.mem[400] [6];
  assign _07612_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [6] : \MSYNC_1r1w.synth.nz.mem[402] [6];
  assign _07613_ = \bapg_rd.w_ptr_r [1] ? _07612_ : _07611_;
  assign _07614_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [6] : \MSYNC_1r1w.synth.nz.mem[404] [6];
  assign _07615_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [6] : \MSYNC_1r1w.synth.nz.mem[406] [6];
  assign _07616_ = \bapg_rd.w_ptr_r [1] ? _07615_ : _07614_;
  assign _07617_ = \bapg_rd.w_ptr_r [2] ? _07616_ : _07613_;
  assign _07618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [6] : \MSYNC_1r1w.synth.nz.mem[408] [6];
  assign _07619_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [6] : \MSYNC_1r1w.synth.nz.mem[410] [6];
  assign _07620_ = \bapg_rd.w_ptr_r [1] ? _07619_ : _07618_;
  assign _07621_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [6] : \MSYNC_1r1w.synth.nz.mem[412] [6];
  assign _07622_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [6] : \MSYNC_1r1w.synth.nz.mem[414] [6];
  assign _07623_ = \bapg_rd.w_ptr_r [1] ? _07622_ : _07621_;
  assign _07624_ = \bapg_rd.w_ptr_r [2] ? _07623_ : _07620_;
  assign _07625_ = \bapg_rd.w_ptr_r [3] ? _07624_ : _07617_;
  assign _07626_ = \bapg_rd.w_ptr_r [4] ? _07625_ : _07610_;
  assign _07627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [6] : \MSYNC_1r1w.synth.nz.mem[416] [6];
  assign _07628_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [6] : \MSYNC_1r1w.synth.nz.mem[418] [6];
  assign _07629_ = \bapg_rd.w_ptr_r [1] ? _07628_ : _07627_;
  assign _07630_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [6] : \MSYNC_1r1w.synth.nz.mem[420] [6];
  assign _07631_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [6] : \MSYNC_1r1w.synth.nz.mem[422] [6];
  assign _07632_ = \bapg_rd.w_ptr_r [1] ? _07631_ : _07630_;
  assign _07633_ = \bapg_rd.w_ptr_r [2] ? _07632_ : _07629_;
  assign _07634_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [6] : \MSYNC_1r1w.synth.nz.mem[424] [6];
  assign _07635_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [6] : \MSYNC_1r1w.synth.nz.mem[426] [6];
  assign _07636_ = \bapg_rd.w_ptr_r [1] ? _07635_ : _07634_;
  assign _07637_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [6] : \MSYNC_1r1w.synth.nz.mem[428] [6];
  assign _07638_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [6] : \MSYNC_1r1w.synth.nz.mem[430] [6];
  assign _07639_ = \bapg_rd.w_ptr_r [1] ? _07638_ : _07637_;
  assign _07640_ = \bapg_rd.w_ptr_r [2] ? _07639_ : _07636_;
  assign _07641_ = \bapg_rd.w_ptr_r [3] ? _07640_ : _07633_;
  assign _07642_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [6] : \MSYNC_1r1w.synth.nz.mem[432] [6];
  assign _07643_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [6] : \MSYNC_1r1w.synth.nz.mem[434] [6];
  assign _07644_ = \bapg_rd.w_ptr_r [1] ? _07643_ : _07642_;
  assign _07645_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [6] : \MSYNC_1r1w.synth.nz.mem[436] [6];
  assign _07646_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [6] : \MSYNC_1r1w.synth.nz.mem[438] [6];
  assign _07647_ = \bapg_rd.w_ptr_r [1] ? _07646_ : _07645_;
  assign _07648_ = \bapg_rd.w_ptr_r [2] ? _07647_ : _07644_;
  assign _07649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [6] : \MSYNC_1r1w.synth.nz.mem[440] [6];
  assign _07650_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [6] : \MSYNC_1r1w.synth.nz.mem[442] [6];
  assign _07651_ = \bapg_rd.w_ptr_r [1] ? _07650_ : _07649_;
  assign _07652_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [6] : \MSYNC_1r1w.synth.nz.mem[444] [6];
  assign _07653_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [6] : \MSYNC_1r1w.synth.nz.mem[446] [6];
  assign _07654_ = \bapg_rd.w_ptr_r [1] ? _07653_ : _07652_;
  assign _07655_ = \bapg_rd.w_ptr_r [2] ? _07654_ : _07651_;
  assign _07656_ = \bapg_rd.w_ptr_r [3] ? _07655_ : _07648_;
  assign _07657_ = \bapg_rd.w_ptr_r [4] ? _07656_ : _07641_;
  assign _07658_ = \bapg_rd.w_ptr_r [5] ? _07657_ : _07626_;
  assign _07659_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [6] : \MSYNC_1r1w.synth.nz.mem[448] [6];
  assign _07660_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [6] : \MSYNC_1r1w.synth.nz.mem[450] [6];
  assign _07661_ = \bapg_rd.w_ptr_r [1] ? _07660_ : _07659_;
  assign _07662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [6] : \MSYNC_1r1w.synth.nz.mem[452] [6];
  assign _07663_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [6] : \MSYNC_1r1w.synth.nz.mem[454] [6];
  assign _07664_ = \bapg_rd.w_ptr_r [1] ? _07663_ : _07662_;
  assign _07665_ = \bapg_rd.w_ptr_r [2] ? _07664_ : _07661_;
  assign _07666_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [6] : \MSYNC_1r1w.synth.nz.mem[456] [6];
  assign _07667_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [6] : \MSYNC_1r1w.synth.nz.mem[458] [6];
  assign _07668_ = \bapg_rd.w_ptr_r [1] ? _07667_ : _07666_;
  assign _07669_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [6] : \MSYNC_1r1w.synth.nz.mem[460] [6];
  assign _07670_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [6] : \MSYNC_1r1w.synth.nz.mem[462] [6];
  assign _07671_ = \bapg_rd.w_ptr_r [1] ? _07670_ : _07669_;
  assign _07672_ = \bapg_rd.w_ptr_r [2] ? _07671_ : _07668_;
  assign _07673_ = \bapg_rd.w_ptr_r [3] ? _07672_ : _07665_;
  assign _07674_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [6] : \MSYNC_1r1w.synth.nz.mem[464] [6];
  assign _07675_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [6] : \MSYNC_1r1w.synth.nz.mem[466] [6];
  assign _07676_ = \bapg_rd.w_ptr_r [1] ? _07675_ : _07674_;
  assign _07677_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [6] : \MSYNC_1r1w.synth.nz.mem[468] [6];
  assign _07678_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [6] : \MSYNC_1r1w.synth.nz.mem[470] [6];
  assign _07679_ = \bapg_rd.w_ptr_r [1] ? _07678_ : _07677_;
  assign _07680_ = \bapg_rd.w_ptr_r [2] ? _07679_ : _07676_;
  assign _07681_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [6] : \MSYNC_1r1w.synth.nz.mem[472] [6];
  assign _07682_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [6] : \MSYNC_1r1w.synth.nz.mem[474] [6];
  assign _07683_ = \bapg_rd.w_ptr_r [1] ? _07682_ : _07681_;
  assign _07684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [6] : \MSYNC_1r1w.synth.nz.mem[476] [6];
  assign _07685_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [6] : \MSYNC_1r1w.synth.nz.mem[478] [6];
  assign _07686_ = \bapg_rd.w_ptr_r [1] ? _07685_ : _07684_;
  assign _07687_ = \bapg_rd.w_ptr_r [2] ? _07686_ : _07683_;
  assign _07688_ = \bapg_rd.w_ptr_r [3] ? _07687_ : _07680_;
  assign _07689_ = \bapg_rd.w_ptr_r [4] ? _07688_ : _07673_;
  assign _07690_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [6] : \MSYNC_1r1w.synth.nz.mem[480] [6];
  assign _07691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [6] : \MSYNC_1r1w.synth.nz.mem[482] [6];
  assign _07692_ = \bapg_rd.w_ptr_r [1] ? _07691_ : _07690_;
  assign _07693_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [6] : \MSYNC_1r1w.synth.nz.mem[484] [6];
  assign _07694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [6] : \MSYNC_1r1w.synth.nz.mem[486] [6];
  assign _07695_ = \bapg_rd.w_ptr_r [1] ? _07694_ : _07693_;
  assign _07696_ = \bapg_rd.w_ptr_r [2] ? _07695_ : _07692_;
  assign _07697_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [6] : \MSYNC_1r1w.synth.nz.mem[488] [6];
  assign _07698_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [6] : \MSYNC_1r1w.synth.nz.mem[490] [6];
  assign _07699_ = \bapg_rd.w_ptr_r [1] ? _07698_ : _07697_;
  assign _07700_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [6] : \MSYNC_1r1w.synth.nz.mem[492] [6];
  assign _07701_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [6] : \MSYNC_1r1w.synth.nz.mem[494] [6];
  assign _07702_ = \bapg_rd.w_ptr_r [1] ? _07701_ : _07700_;
  assign _07703_ = \bapg_rd.w_ptr_r [2] ? _07702_ : _07699_;
  assign _07704_ = \bapg_rd.w_ptr_r [3] ? _07703_ : _07696_;
  assign _07705_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [6] : \MSYNC_1r1w.synth.nz.mem[496] [6];
  assign _07706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [6] : \MSYNC_1r1w.synth.nz.mem[498] [6];
  assign _07707_ = \bapg_rd.w_ptr_r [1] ? _07706_ : _07705_;
  assign _07708_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [6] : \MSYNC_1r1w.synth.nz.mem[500] [6];
  assign _07709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [6] : \MSYNC_1r1w.synth.nz.mem[502] [6];
  assign _07710_ = \bapg_rd.w_ptr_r [1] ? _07709_ : _07708_;
  assign _07711_ = \bapg_rd.w_ptr_r [2] ? _07710_ : _07707_;
  assign _07712_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [6] : \MSYNC_1r1w.synth.nz.mem[504] [6];
  assign _07713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [6] : \MSYNC_1r1w.synth.nz.mem[506] [6];
  assign _07714_ = \bapg_rd.w_ptr_r [1] ? _07713_ : _07712_;
  assign _07715_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [6] : \MSYNC_1r1w.synth.nz.mem[508] [6];
  assign _07716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [6] : \MSYNC_1r1w.synth.nz.mem[510] [6];
  assign _07717_ = \bapg_rd.w_ptr_r [1] ? _07716_ : _07715_;
  assign _07718_ = \bapg_rd.w_ptr_r [2] ? _07717_ : _07714_;
  assign _07719_ = \bapg_rd.w_ptr_r [3] ? _07718_ : _07711_;
  assign _07720_ = \bapg_rd.w_ptr_r [4] ? _07719_ : _07704_;
  assign _07721_ = \bapg_rd.w_ptr_r [5] ? _07720_ : _07689_;
  assign _07722_ = \bapg_rd.w_ptr_r [6] ? _07721_ : _07658_;
  assign _07723_ = \bapg_rd.w_ptr_r [7] ? _07722_ : _07595_;
  assign _07724_ = \bapg_rd.w_ptr_r [8] ? _07723_ : _07468_;
  assign _07725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [6] : \MSYNC_1r1w.synth.nz.mem[512] [6];
  assign _07726_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [6] : \MSYNC_1r1w.synth.nz.mem[514] [6];
  assign _07727_ = \bapg_rd.w_ptr_r [1] ? _07726_ : _07725_;
  assign _07728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [6] : \MSYNC_1r1w.synth.nz.mem[516] [6];
  assign _07729_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [6] : \MSYNC_1r1w.synth.nz.mem[518] [6];
  assign _07730_ = \bapg_rd.w_ptr_r [1] ? _07729_ : _07728_;
  assign _07731_ = \bapg_rd.w_ptr_r [2] ? _07730_ : _07727_;
  assign _07732_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [6] : \MSYNC_1r1w.synth.nz.mem[520] [6];
  assign _07733_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [6] : \MSYNC_1r1w.synth.nz.mem[522] [6];
  assign _07734_ = \bapg_rd.w_ptr_r [1] ? _07733_ : _07732_;
  assign _07735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [6] : \MSYNC_1r1w.synth.nz.mem[524] [6];
  assign _07736_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [6] : \MSYNC_1r1w.synth.nz.mem[526] [6];
  assign _07737_ = \bapg_rd.w_ptr_r [1] ? _07736_ : _07735_;
  assign _07738_ = \bapg_rd.w_ptr_r [2] ? _07737_ : _07734_;
  assign _07739_ = \bapg_rd.w_ptr_r [3] ? _07738_ : _07731_;
  assign _07740_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [6] : \MSYNC_1r1w.synth.nz.mem[528] [6];
  assign _07741_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [6] : \MSYNC_1r1w.synth.nz.mem[530] [6];
  assign _07742_ = \bapg_rd.w_ptr_r [1] ? _07741_ : _07740_;
  assign _07743_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [6] : \MSYNC_1r1w.synth.nz.mem[532] [6];
  assign _07744_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [6] : \MSYNC_1r1w.synth.nz.mem[534] [6];
  assign _07745_ = \bapg_rd.w_ptr_r [1] ? _07744_ : _07743_;
  assign _07746_ = \bapg_rd.w_ptr_r [2] ? _07745_ : _07742_;
  assign _07747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [6] : \MSYNC_1r1w.synth.nz.mem[536] [6];
  assign _07748_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [6] : \MSYNC_1r1w.synth.nz.mem[538] [6];
  assign _07749_ = \bapg_rd.w_ptr_r [1] ? _07748_ : _07747_;
  assign _07750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [6] : \MSYNC_1r1w.synth.nz.mem[540] [6];
  assign _07751_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [6] : \MSYNC_1r1w.synth.nz.mem[542] [6];
  assign _07752_ = \bapg_rd.w_ptr_r [1] ? _07751_ : _07750_;
  assign _07753_ = \bapg_rd.w_ptr_r [2] ? _07752_ : _07749_;
  assign _07754_ = \bapg_rd.w_ptr_r [3] ? _07753_ : _07746_;
  assign _07755_ = \bapg_rd.w_ptr_r [4] ? _07754_ : _07739_;
  assign _07756_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [6] : \MSYNC_1r1w.synth.nz.mem[544] [6];
  assign _07757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [6] : \MSYNC_1r1w.synth.nz.mem[546] [6];
  assign _07758_ = \bapg_rd.w_ptr_r [1] ? _07757_ : _07756_;
  assign _07759_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [6] : \MSYNC_1r1w.synth.nz.mem[548] [6];
  assign _07760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [6] : \MSYNC_1r1w.synth.nz.mem[550] [6];
  assign _07761_ = \bapg_rd.w_ptr_r [1] ? _07760_ : _07759_;
  assign _07762_ = \bapg_rd.w_ptr_r [2] ? _07761_ : _07758_;
  assign _07763_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [6] : \MSYNC_1r1w.synth.nz.mem[552] [6];
  assign _07764_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [6] : \MSYNC_1r1w.synth.nz.mem[554] [6];
  assign _07765_ = \bapg_rd.w_ptr_r [1] ? _07764_ : _07763_;
  assign _07766_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [6] : \MSYNC_1r1w.synth.nz.mem[556] [6];
  assign _07767_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [6] : \MSYNC_1r1w.synth.nz.mem[558] [6];
  assign _07768_ = \bapg_rd.w_ptr_r [1] ? _07767_ : _07766_;
  assign _07769_ = \bapg_rd.w_ptr_r [2] ? _07768_ : _07765_;
  assign _07770_ = \bapg_rd.w_ptr_r [3] ? _07769_ : _07762_;
  assign _07771_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [6] : \MSYNC_1r1w.synth.nz.mem[560] [6];
  assign _07772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [6] : \MSYNC_1r1w.synth.nz.mem[562] [6];
  assign _07773_ = \bapg_rd.w_ptr_r [1] ? _07772_ : _07771_;
  assign _07774_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [6] : \MSYNC_1r1w.synth.nz.mem[564] [6];
  assign _07775_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [6] : \MSYNC_1r1w.synth.nz.mem[566] [6];
  assign _07776_ = \bapg_rd.w_ptr_r [1] ? _07775_ : _07774_;
  assign _07777_ = \bapg_rd.w_ptr_r [2] ? _07776_ : _07773_;
  assign _07778_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [6] : \MSYNC_1r1w.synth.nz.mem[568] [6];
  assign _07779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [6] : \MSYNC_1r1w.synth.nz.mem[570] [6];
  assign _07780_ = \bapg_rd.w_ptr_r [1] ? _07779_ : _07778_;
  assign _07781_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [6] : \MSYNC_1r1w.synth.nz.mem[572] [6];
  assign _07782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [6] : \MSYNC_1r1w.synth.nz.mem[574] [6];
  assign _07783_ = \bapg_rd.w_ptr_r [1] ? _07782_ : _07781_;
  assign _07784_ = \bapg_rd.w_ptr_r [2] ? _07783_ : _07780_;
  assign _07785_ = \bapg_rd.w_ptr_r [3] ? _07784_ : _07777_;
  assign _07786_ = \bapg_rd.w_ptr_r [4] ? _07785_ : _07770_;
  assign _07787_ = \bapg_rd.w_ptr_r [5] ? _07786_ : _07755_;
  assign _07788_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [6] : \MSYNC_1r1w.synth.nz.mem[576] [6];
  assign _07789_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [6] : \MSYNC_1r1w.synth.nz.mem[578] [6];
  assign _07790_ = \bapg_rd.w_ptr_r [1] ? _07789_ : _07788_;
  assign _07791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [6] : \MSYNC_1r1w.synth.nz.mem[580] [6];
  assign _07792_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [6] : \MSYNC_1r1w.synth.nz.mem[582] [6];
  assign _07793_ = \bapg_rd.w_ptr_r [1] ? _07792_ : _07791_;
  assign _07794_ = \bapg_rd.w_ptr_r [2] ? _07793_ : _07790_;
  assign _07795_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [6] : \MSYNC_1r1w.synth.nz.mem[584] [6];
  assign _07796_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [6] : \MSYNC_1r1w.synth.nz.mem[586] [6];
  assign _07797_ = \bapg_rd.w_ptr_r [1] ? _07796_ : _07795_;
  assign _07798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [6] : \MSYNC_1r1w.synth.nz.mem[588] [6];
  assign _07799_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [6] : \MSYNC_1r1w.synth.nz.mem[590] [6];
  assign _07800_ = \bapg_rd.w_ptr_r [1] ? _07799_ : _07798_;
  assign _07801_ = \bapg_rd.w_ptr_r [2] ? _07800_ : _07797_;
  assign _07802_ = \bapg_rd.w_ptr_r [3] ? _07801_ : _07794_;
  assign _07803_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [6] : \MSYNC_1r1w.synth.nz.mem[592] [6];
  assign _07804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [6] : \MSYNC_1r1w.synth.nz.mem[594] [6];
  assign _07805_ = \bapg_rd.w_ptr_r [1] ? _07804_ : _07803_;
  assign _07806_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [6] : \MSYNC_1r1w.synth.nz.mem[596] [6];
  assign _07807_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [6] : \MSYNC_1r1w.synth.nz.mem[598] [6];
  assign _07808_ = \bapg_rd.w_ptr_r [1] ? _07807_ : _07806_;
  assign _07809_ = \bapg_rd.w_ptr_r [2] ? _07808_ : _07805_;
  assign _07810_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [6] : \MSYNC_1r1w.synth.nz.mem[600] [6];
  assign _07811_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [6] : \MSYNC_1r1w.synth.nz.mem[602] [6];
  assign _07812_ = \bapg_rd.w_ptr_r [1] ? _07811_ : _07810_;
  assign _07813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [6] : \MSYNC_1r1w.synth.nz.mem[604] [6];
  assign _07814_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [6] : \MSYNC_1r1w.synth.nz.mem[606] [6];
  assign _07815_ = \bapg_rd.w_ptr_r [1] ? _07814_ : _07813_;
  assign _07816_ = \bapg_rd.w_ptr_r [2] ? _07815_ : _07812_;
  assign _07817_ = \bapg_rd.w_ptr_r [3] ? _07816_ : _07809_;
  assign _07818_ = \bapg_rd.w_ptr_r [4] ? _07817_ : _07802_;
  assign _07819_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [6] : \MSYNC_1r1w.synth.nz.mem[608] [6];
  assign _07820_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [6] : \MSYNC_1r1w.synth.nz.mem[610] [6];
  assign _07821_ = \bapg_rd.w_ptr_r [1] ? _07820_ : _07819_;
  assign _07822_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [6] : \MSYNC_1r1w.synth.nz.mem[612] [6];
  assign _07823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [6] : \MSYNC_1r1w.synth.nz.mem[614] [6];
  assign _07824_ = \bapg_rd.w_ptr_r [1] ? _07823_ : _07822_;
  assign _07825_ = \bapg_rd.w_ptr_r [2] ? _07824_ : _07821_;
  assign _07826_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [6] : \MSYNC_1r1w.synth.nz.mem[616] [6];
  assign _07827_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [6] : \MSYNC_1r1w.synth.nz.mem[618] [6];
  assign _07828_ = \bapg_rd.w_ptr_r [1] ? _07827_ : _07826_;
  assign _07829_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [6] : \MSYNC_1r1w.synth.nz.mem[620] [6];
  assign _07830_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [6] : \MSYNC_1r1w.synth.nz.mem[622] [6];
  assign _07831_ = \bapg_rd.w_ptr_r [1] ? _07830_ : _07829_;
  assign _07832_ = \bapg_rd.w_ptr_r [2] ? _07831_ : _07828_;
  assign _07833_ = \bapg_rd.w_ptr_r [3] ? _07832_ : _07825_;
  assign _07834_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [6] : \MSYNC_1r1w.synth.nz.mem[624] [6];
  assign _07835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [6] : \MSYNC_1r1w.synth.nz.mem[626] [6];
  assign _07836_ = \bapg_rd.w_ptr_r [1] ? _07835_ : _07834_;
  assign _07837_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [6] : \MSYNC_1r1w.synth.nz.mem[628] [6];
  assign _07838_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [6] : \MSYNC_1r1w.synth.nz.mem[630] [6];
  assign _07839_ = \bapg_rd.w_ptr_r [1] ? _07838_ : _07837_;
  assign _07840_ = \bapg_rd.w_ptr_r [2] ? _07839_ : _07836_;
  assign _07841_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [6] : \MSYNC_1r1w.synth.nz.mem[632] [6];
  assign _07842_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [6] : \MSYNC_1r1w.synth.nz.mem[634] [6];
  assign _07843_ = \bapg_rd.w_ptr_r [1] ? _07842_ : _07841_;
  assign _07844_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [6] : \MSYNC_1r1w.synth.nz.mem[636] [6];
  assign _07845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [6] : \MSYNC_1r1w.synth.nz.mem[638] [6];
  assign _07846_ = \bapg_rd.w_ptr_r [1] ? _07845_ : _07844_;
  assign _07847_ = \bapg_rd.w_ptr_r [2] ? _07846_ : _07843_;
  assign _07848_ = \bapg_rd.w_ptr_r [3] ? _07847_ : _07840_;
  assign _07849_ = \bapg_rd.w_ptr_r [4] ? _07848_ : _07833_;
  assign _07850_ = \bapg_rd.w_ptr_r [5] ? _07849_ : _07818_;
  assign _07851_ = \bapg_rd.w_ptr_r [6] ? _07850_ : _07787_;
  assign _07852_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [6] : \MSYNC_1r1w.synth.nz.mem[640] [6];
  assign _07853_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [6] : \MSYNC_1r1w.synth.nz.mem[642] [6];
  assign _07854_ = \bapg_rd.w_ptr_r [1] ? _07853_ : _07852_;
  assign _07855_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [6] : \MSYNC_1r1w.synth.nz.mem[644] [6];
  assign _07856_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [6] : \MSYNC_1r1w.synth.nz.mem[646] [6];
  assign _07857_ = \bapg_rd.w_ptr_r [1] ? _07856_ : _07855_;
  assign _07858_ = \bapg_rd.w_ptr_r [2] ? _07857_ : _07854_;
  assign _07859_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [6] : \MSYNC_1r1w.synth.nz.mem[648] [6];
  assign _07860_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [6] : \MSYNC_1r1w.synth.nz.mem[650] [6];
  assign _07861_ = \bapg_rd.w_ptr_r [1] ? _07860_ : _07859_;
  assign _07862_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [6] : \MSYNC_1r1w.synth.nz.mem[652] [6];
  assign _07863_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [6] : \MSYNC_1r1w.synth.nz.mem[654] [6];
  assign _07864_ = \bapg_rd.w_ptr_r [1] ? _07863_ : _07862_;
  assign _07865_ = \bapg_rd.w_ptr_r [2] ? _07864_ : _07861_;
  assign _07866_ = \bapg_rd.w_ptr_r [3] ? _07865_ : _07858_;
  assign _07867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [6] : \MSYNC_1r1w.synth.nz.mem[656] [6];
  assign _07868_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [6] : \MSYNC_1r1w.synth.nz.mem[658] [6];
  assign _07869_ = \bapg_rd.w_ptr_r [1] ? _07868_ : _07867_;
  assign _07870_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [6] : \MSYNC_1r1w.synth.nz.mem[660] [6];
  assign _07871_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [6] : \MSYNC_1r1w.synth.nz.mem[662] [6];
  assign _07872_ = \bapg_rd.w_ptr_r [1] ? _07871_ : _07870_;
  assign _07873_ = \bapg_rd.w_ptr_r [2] ? _07872_ : _07869_;
  assign _07874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [6] : \MSYNC_1r1w.synth.nz.mem[664] [6];
  assign _07875_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [6] : \MSYNC_1r1w.synth.nz.mem[666] [6];
  assign _07876_ = \bapg_rd.w_ptr_r [1] ? _07875_ : _07874_;
  assign _07877_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [6] : \MSYNC_1r1w.synth.nz.mem[668] [6];
  assign _07878_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [6] : \MSYNC_1r1w.synth.nz.mem[670] [6];
  assign _07879_ = \bapg_rd.w_ptr_r [1] ? _07878_ : _07877_;
  assign _07880_ = \bapg_rd.w_ptr_r [2] ? _07879_ : _07876_;
  assign _07881_ = \bapg_rd.w_ptr_r [3] ? _07880_ : _07873_;
  assign _07882_ = \bapg_rd.w_ptr_r [4] ? _07881_ : _07866_;
  assign _07883_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [6] : \MSYNC_1r1w.synth.nz.mem[672] [6];
  assign _07884_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [6] : \MSYNC_1r1w.synth.nz.mem[674] [6];
  assign _07885_ = \bapg_rd.w_ptr_r [1] ? _07884_ : _07883_;
  assign _07886_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [6] : \MSYNC_1r1w.synth.nz.mem[676] [6];
  assign _07887_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [6] : \MSYNC_1r1w.synth.nz.mem[678] [6];
  assign _07888_ = \bapg_rd.w_ptr_r [1] ? _07887_ : _07886_;
  assign _07889_ = \bapg_rd.w_ptr_r [2] ? _07888_ : _07885_;
  assign _07890_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [6] : \MSYNC_1r1w.synth.nz.mem[680] [6];
  assign _07891_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [6] : \MSYNC_1r1w.synth.nz.mem[682] [6];
  assign _07892_ = \bapg_rd.w_ptr_r [1] ? _07891_ : _07890_;
  assign _07893_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [6] : \MSYNC_1r1w.synth.nz.mem[684] [6];
  assign _07894_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [6] : \MSYNC_1r1w.synth.nz.mem[686] [6];
  assign _07895_ = \bapg_rd.w_ptr_r [1] ? _07894_ : _07893_;
  assign _07896_ = \bapg_rd.w_ptr_r [2] ? _07895_ : _07892_;
  assign _07897_ = \bapg_rd.w_ptr_r [3] ? _07896_ : _07889_;
  assign _07898_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [6] : \MSYNC_1r1w.synth.nz.mem[688] [6];
  assign _07899_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [6] : \MSYNC_1r1w.synth.nz.mem[690] [6];
  assign _07900_ = \bapg_rd.w_ptr_r [1] ? _07899_ : _07898_;
  assign _07901_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [6] : \MSYNC_1r1w.synth.nz.mem[692] [6];
  assign _07902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [6] : \MSYNC_1r1w.synth.nz.mem[694] [6];
  assign _07903_ = \bapg_rd.w_ptr_r [1] ? _07902_ : _07901_;
  assign _07904_ = \bapg_rd.w_ptr_r [2] ? _07903_ : _07900_;
  assign _07905_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [6] : \MSYNC_1r1w.synth.nz.mem[696] [6];
  assign _07906_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [6] : \MSYNC_1r1w.synth.nz.mem[698] [6];
  assign _07907_ = \bapg_rd.w_ptr_r [1] ? _07906_ : _07905_;
  assign _07908_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [6] : \MSYNC_1r1w.synth.nz.mem[700] [6];
  assign _07909_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [6] : \MSYNC_1r1w.synth.nz.mem[702] [6];
  assign _07910_ = \bapg_rd.w_ptr_r [1] ? _07909_ : _07908_;
  assign _07911_ = \bapg_rd.w_ptr_r [2] ? _07910_ : _07907_;
  assign _07912_ = \bapg_rd.w_ptr_r [3] ? _07911_ : _07904_;
  assign _07913_ = \bapg_rd.w_ptr_r [4] ? _07912_ : _07897_;
  assign _07914_ = \bapg_rd.w_ptr_r [5] ? _07913_ : _07882_;
  assign _07915_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [6] : \MSYNC_1r1w.synth.nz.mem[704] [6];
  assign _07916_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [6] : \MSYNC_1r1w.synth.nz.mem[706] [6];
  assign _07917_ = \bapg_rd.w_ptr_r [1] ? _07916_ : _07915_;
  assign _07918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [6] : \MSYNC_1r1w.synth.nz.mem[708] [6];
  assign _07919_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [6] : \MSYNC_1r1w.synth.nz.mem[710] [6];
  assign _07920_ = \bapg_rd.w_ptr_r [1] ? _07919_ : _07918_;
  assign _07921_ = \bapg_rd.w_ptr_r [2] ? _07920_ : _07917_;
  assign _07922_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [6] : \MSYNC_1r1w.synth.nz.mem[712] [6];
  assign _07923_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [6] : \MSYNC_1r1w.synth.nz.mem[714] [6];
  assign _07924_ = \bapg_rd.w_ptr_r [1] ? _07923_ : _07922_;
  assign _07925_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [6] : \MSYNC_1r1w.synth.nz.mem[716] [6];
  assign _07926_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [6] : \MSYNC_1r1w.synth.nz.mem[718] [6];
  assign _07927_ = \bapg_rd.w_ptr_r [1] ? _07926_ : _07925_;
  assign _07928_ = \bapg_rd.w_ptr_r [2] ? _07927_ : _07924_;
  assign _07929_ = \bapg_rd.w_ptr_r [3] ? _07928_ : _07921_;
  assign _07930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [6] : \MSYNC_1r1w.synth.nz.mem[720] [6];
  assign _07931_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [6] : \MSYNC_1r1w.synth.nz.mem[722] [6];
  assign _07932_ = \bapg_rd.w_ptr_r [1] ? _07931_ : _07930_;
  assign _07933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [6] : \MSYNC_1r1w.synth.nz.mem[724] [6];
  assign _07934_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [6] : \MSYNC_1r1w.synth.nz.mem[726] [6];
  assign _07935_ = \bapg_rd.w_ptr_r [1] ? _07934_ : _07933_;
  assign _07936_ = \bapg_rd.w_ptr_r [2] ? _07935_ : _07932_;
  assign _07937_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [6] : \MSYNC_1r1w.synth.nz.mem[728] [6];
  assign _07938_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [6] : \MSYNC_1r1w.synth.nz.mem[730] [6];
  assign _07939_ = \bapg_rd.w_ptr_r [1] ? _07938_ : _07937_;
  assign _07940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [6] : \MSYNC_1r1w.synth.nz.mem[732] [6];
  assign _07941_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [6] : \MSYNC_1r1w.synth.nz.mem[734] [6];
  assign _07942_ = \bapg_rd.w_ptr_r [1] ? _07941_ : _07940_;
  assign _07943_ = \bapg_rd.w_ptr_r [2] ? _07942_ : _07939_;
  assign _07944_ = \bapg_rd.w_ptr_r [3] ? _07943_ : _07936_;
  assign _07945_ = \bapg_rd.w_ptr_r [4] ? _07944_ : _07929_;
  assign _07946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [6] : \MSYNC_1r1w.synth.nz.mem[736] [6];
  assign _07947_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [6] : \MSYNC_1r1w.synth.nz.mem[738] [6];
  assign _07948_ = \bapg_rd.w_ptr_r [1] ? _07947_ : _07946_;
  assign _07949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [6] : \MSYNC_1r1w.synth.nz.mem[740] [6];
  assign _07950_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [6] : \MSYNC_1r1w.synth.nz.mem[742] [6];
  assign _07951_ = \bapg_rd.w_ptr_r [1] ? _07950_ : _07949_;
  assign _07952_ = \bapg_rd.w_ptr_r [2] ? _07951_ : _07948_;
  assign _07953_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [6] : \MSYNC_1r1w.synth.nz.mem[744] [6];
  assign _07954_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [6] : \MSYNC_1r1w.synth.nz.mem[746] [6];
  assign _07955_ = \bapg_rd.w_ptr_r [1] ? _07954_ : _07953_;
  assign _07956_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [6] : \MSYNC_1r1w.synth.nz.mem[748] [6];
  assign _07957_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [6] : \MSYNC_1r1w.synth.nz.mem[750] [6];
  assign _07958_ = \bapg_rd.w_ptr_r [1] ? _07957_ : _07956_;
  assign _07959_ = \bapg_rd.w_ptr_r [2] ? _07958_ : _07955_;
  assign _07960_ = \bapg_rd.w_ptr_r [3] ? _07959_ : _07952_;
  assign _07961_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [6] : \MSYNC_1r1w.synth.nz.mem[752] [6];
  assign _07962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [6] : \MSYNC_1r1w.synth.nz.mem[754] [6];
  assign _07963_ = \bapg_rd.w_ptr_r [1] ? _07962_ : _07961_;
  assign _07964_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [6] : \MSYNC_1r1w.synth.nz.mem[756] [6];
  assign _07965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [6] : \MSYNC_1r1w.synth.nz.mem[758] [6];
  assign _07966_ = \bapg_rd.w_ptr_r [1] ? _07965_ : _07964_;
  assign _07967_ = \bapg_rd.w_ptr_r [2] ? _07966_ : _07963_;
  assign _07968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [6] : \MSYNC_1r1w.synth.nz.mem[760] [6];
  assign _07969_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [6] : \MSYNC_1r1w.synth.nz.mem[762] [6];
  assign _07970_ = \bapg_rd.w_ptr_r [1] ? _07969_ : _07968_;
  assign _07971_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [6] : \MSYNC_1r1w.synth.nz.mem[764] [6];
  assign _07972_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [6] : \MSYNC_1r1w.synth.nz.mem[766] [6];
  assign _07973_ = \bapg_rd.w_ptr_r [1] ? _07972_ : _07971_;
  assign _07974_ = \bapg_rd.w_ptr_r [2] ? _07973_ : _07970_;
  assign _07975_ = \bapg_rd.w_ptr_r [3] ? _07974_ : _07967_;
  assign _07976_ = \bapg_rd.w_ptr_r [4] ? _07975_ : _07960_;
  assign _07977_ = \bapg_rd.w_ptr_r [5] ? _07976_ : _07945_;
  assign _07978_ = \bapg_rd.w_ptr_r [6] ? _07977_ : _07914_;
  assign _07979_ = \bapg_rd.w_ptr_r [7] ? _07978_ : _07851_;
  assign _07980_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [6] : \MSYNC_1r1w.synth.nz.mem[768] [6];
  assign _07981_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [6] : \MSYNC_1r1w.synth.nz.mem[770] [6];
  assign _07982_ = \bapg_rd.w_ptr_r [1] ? _07981_ : _07980_;
  assign _07983_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [6] : \MSYNC_1r1w.synth.nz.mem[772] [6];
  assign _07984_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [6] : \MSYNC_1r1w.synth.nz.mem[774] [6];
  assign _07985_ = \bapg_rd.w_ptr_r [1] ? _07984_ : _07983_;
  assign _07986_ = \bapg_rd.w_ptr_r [2] ? _07985_ : _07982_;
  assign _07987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [6] : \MSYNC_1r1w.synth.nz.mem[776] [6];
  assign _07988_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [6] : \MSYNC_1r1w.synth.nz.mem[778] [6];
  assign _07989_ = \bapg_rd.w_ptr_r [1] ? _07988_ : _07987_;
  assign _07990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [6] : \MSYNC_1r1w.synth.nz.mem[780] [6];
  assign _07991_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [6] : \MSYNC_1r1w.synth.nz.mem[782] [6];
  assign _07992_ = \bapg_rd.w_ptr_r [1] ? _07991_ : _07990_;
  assign _07993_ = \bapg_rd.w_ptr_r [2] ? _07992_ : _07989_;
  assign _07994_ = \bapg_rd.w_ptr_r [3] ? _07993_ : _07986_;
  assign _07995_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [6] : \MSYNC_1r1w.synth.nz.mem[784] [6];
  assign _07996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [6] : \MSYNC_1r1w.synth.nz.mem[786] [6];
  assign _07997_ = \bapg_rd.w_ptr_r [1] ? _07996_ : _07995_;
  assign _07998_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [6] : \MSYNC_1r1w.synth.nz.mem[788] [6];
  assign _07999_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [6] : \MSYNC_1r1w.synth.nz.mem[790] [6];
  assign _08000_ = \bapg_rd.w_ptr_r [1] ? _07999_ : _07998_;
  assign _08001_ = \bapg_rd.w_ptr_r [2] ? _08000_ : _07997_;
  assign _08002_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [6] : \MSYNC_1r1w.synth.nz.mem[792] [6];
  assign _08003_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [6] : \MSYNC_1r1w.synth.nz.mem[794] [6];
  assign _08004_ = \bapg_rd.w_ptr_r [1] ? _08003_ : _08002_;
  assign _08005_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [6] : \MSYNC_1r1w.synth.nz.mem[796] [6];
  assign _08006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [6] : \MSYNC_1r1w.synth.nz.mem[798] [6];
  assign _08007_ = \bapg_rd.w_ptr_r [1] ? _08006_ : _08005_;
  assign _08008_ = \bapg_rd.w_ptr_r [2] ? _08007_ : _08004_;
  assign _08009_ = \bapg_rd.w_ptr_r [3] ? _08008_ : _08001_;
  assign _08010_ = \bapg_rd.w_ptr_r [4] ? _08009_ : _07994_;
  assign _08011_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [6] : \MSYNC_1r1w.synth.nz.mem[800] [6];
  assign _08012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [6] : \MSYNC_1r1w.synth.nz.mem[802] [6];
  assign _08013_ = \bapg_rd.w_ptr_r [1] ? _08012_ : _08011_;
  assign _08014_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [6] : \MSYNC_1r1w.synth.nz.mem[804] [6];
  assign _08015_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [6] : \MSYNC_1r1w.synth.nz.mem[806] [6];
  assign _08016_ = \bapg_rd.w_ptr_r [1] ? _08015_ : _08014_;
  assign _08017_ = \bapg_rd.w_ptr_r [2] ? _08016_ : _08013_;
  assign _08018_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [6] : \MSYNC_1r1w.synth.nz.mem[808] [6];
  assign _08019_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [6] : \MSYNC_1r1w.synth.nz.mem[810] [6];
  assign _08020_ = \bapg_rd.w_ptr_r [1] ? _08019_ : _08018_;
  assign _08021_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [6] : \MSYNC_1r1w.synth.nz.mem[812] [6];
  assign _08022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [6] : \MSYNC_1r1w.synth.nz.mem[814] [6];
  assign _08023_ = \bapg_rd.w_ptr_r [1] ? _08022_ : _08021_;
  assign _08024_ = \bapg_rd.w_ptr_r [2] ? _08023_ : _08020_;
  assign _08025_ = \bapg_rd.w_ptr_r [3] ? _08024_ : _08017_;
  assign _08026_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [6] : \MSYNC_1r1w.synth.nz.mem[816] [6];
  assign _08027_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [6] : \MSYNC_1r1w.synth.nz.mem[818] [6];
  assign _08028_ = \bapg_rd.w_ptr_r [1] ? _08027_ : _08026_;
  assign _08029_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [6] : \MSYNC_1r1w.synth.nz.mem[820] [6];
  assign _08030_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [6] : \MSYNC_1r1w.synth.nz.mem[822] [6];
  assign _08031_ = \bapg_rd.w_ptr_r [1] ? _08030_ : _08029_;
  assign _08032_ = \bapg_rd.w_ptr_r [2] ? _08031_ : _08028_;
  assign _08033_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [6] : \MSYNC_1r1w.synth.nz.mem[824] [6];
  assign _08034_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [6] : \MSYNC_1r1w.synth.nz.mem[826] [6];
  assign _08035_ = \bapg_rd.w_ptr_r [1] ? _08034_ : _08033_;
  assign _08036_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [6] : \MSYNC_1r1w.synth.nz.mem[828] [6];
  assign _08037_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [6] : \MSYNC_1r1w.synth.nz.mem[830] [6];
  assign _08038_ = \bapg_rd.w_ptr_r [1] ? _08037_ : _08036_;
  assign _08039_ = \bapg_rd.w_ptr_r [2] ? _08038_ : _08035_;
  assign _08040_ = \bapg_rd.w_ptr_r [3] ? _08039_ : _08032_;
  assign _08041_ = \bapg_rd.w_ptr_r [4] ? _08040_ : _08025_;
  assign _08042_ = \bapg_rd.w_ptr_r [5] ? _08041_ : _08010_;
  assign _08043_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [6] : \MSYNC_1r1w.synth.nz.mem[832] [6];
  assign _08044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [6] : \MSYNC_1r1w.synth.nz.mem[834] [6];
  assign _08045_ = \bapg_rd.w_ptr_r [1] ? _08044_ : _08043_;
  assign _08046_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [6] : \MSYNC_1r1w.synth.nz.mem[836] [6];
  assign _08047_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [6] : \MSYNC_1r1w.synth.nz.mem[838] [6];
  assign _08048_ = \bapg_rd.w_ptr_r [1] ? _08047_ : _08046_;
  assign _08049_ = \bapg_rd.w_ptr_r [2] ? _08048_ : _08045_;
  assign _08050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [6] : \MSYNC_1r1w.synth.nz.mem[840] [6];
  assign _08051_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [6] : \MSYNC_1r1w.synth.nz.mem[842] [6];
  assign _08052_ = \bapg_rd.w_ptr_r [1] ? _08051_ : _08050_;
  assign _08053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [6] : \MSYNC_1r1w.synth.nz.mem[844] [6];
  assign _08054_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [6] : \MSYNC_1r1w.synth.nz.mem[846] [6];
  assign _08055_ = \bapg_rd.w_ptr_r [1] ? _08054_ : _08053_;
  assign _08056_ = \bapg_rd.w_ptr_r [2] ? _08055_ : _08052_;
  assign _08057_ = \bapg_rd.w_ptr_r [3] ? _08056_ : _08049_;
  assign _08058_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [6] : \MSYNC_1r1w.synth.nz.mem[848] [6];
  assign _08059_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [6] : \MSYNC_1r1w.synth.nz.mem[850] [6];
  assign _08060_ = \bapg_rd.w_ptr_r [1] ? _08059_ : _08058_;
  assign _08061_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [6] : \MSYNC_1r1w.synth.nz.mem[852] [6];
  assign _08062_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [6] : \MSYNC_1r1w.synth.nz.mem[854] [6];
  assign _08063_ = \bapg_rd.w_ptr_r [1] ? _08062_ : _08061_;
  assign _08064_ = \bapg_rd.w_ptr_r [2] ? _08063_ : _08060_;
  assign _08065_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [6] : \MSYNC_1r1w.synth.nz.mem[856] [6];
  assign _08066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [6] : \MSYNC_1r1w.synth.nz.mem[858] [6];
  assign _08067_ = \bapg_rd.w_ptr_r [1] ? _08066_ : _08065_;
  assign _08068_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [6] : \MSYNC_1r1w.synth.nz.mem[860] [6];
  assign _08069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [6] : \MSYNC_1r1w.synth.nz.mem[862] [6];
  assign _08070_ = \bapg_rd.w_ptr_r [1] ? _08069_ : _08068_;
  assign _08071_ = \bapg_rd.w_ptr_r [2] ? _08070_ : _08067_;
  assign _08072_ = \bapg_rd.w_ptr_r [3] ? _08071_ : _08064_;
  assign _08073_ = \bapg_rd.w_ptr_r [4] ? _08072_ : _08057_;
  assign _08074_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [6] : \MSYNC_1r1w.synth.nz.mem[864] [6];
  assign _08075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [6] : \MSYNC_1r1w.synth.nz.mem[866] [6];
  assign _08076_ = \bapg_rd.w_ptr_r [1] ? _08075_ : _08074_;
  assign _08077_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [6] : \MSYNC_1r1w.synth.nz.mem[868] [6];
  assign _08078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [6] : \MSYNC_1r1w.synth.nz.mem[870] [6];
  assign _08079_ = \bapg_rd.w_ptr_r [1] ? _08078_ : _08077_;
  assign _08080_ = \bapg_rd.w_ptr_r [2] ? _08079_ : _08076_;
  assign _08081_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [6] : \MSYNC_1r1w.synth.nz.mem[872] [6];
  assign _08082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [6] : \MSYNC_1r1w.synth.nz.mem[874] [6];
  assign _08083_ = \bapg_rd.w_ptr_r [1] ? _08082_ : _08081_;
  assign _08084_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [6] : \MSYNC_1r1w.synth.nz.mem[876] [6];
  assign _08085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [6] : \MSYNC_1r1w.synth.nz.mem[878] [6];
  assign _08086_ = \bapg_rd.w_ptr_r [1] ? _08085_ : _08084_;
  assign _08087_ = \bapg_rd.w_ptr_r [2] ? _08086_ : _08083_;
  assign _08088_ = \bapg_rd.w_ptr_r [3] ? _08087_ : _08080_;
  assign _08089_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [6] : \MSYNC_1r1w.synth.nz.mem[880] [6];
  assign _08090_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [6] : \MSYNC_1r1w.synth.nz.mem[882] [6];
  assign _08091_ = \bapg_rd.w_ptr_r [1] ? _08090_ : _08089_;
  assign _08092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [6] : \MSYNC_1r1w.synth.nz.mem[884] [6];
  assign _08093_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [6] : \MSYNC_1r1w.synth.nz.mem[886] [6];
  assign _08094_ = \bapg_rd.w_ptr_r [1] ? _08093_ : _08092_;
  assign _08095_ = \bapg_rd.w_ptr_r [2] ? _08094_ : _08091_;
  assign _08096_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [6] : \MSYNC_1r1w.synth.nz.mem[888] [6];
  assign _08097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [6] : \MSYNC_1r1w.synth.nz.mem[890] [6];
  assign _08098_ = \bapg_rd.w_ptr_r [1] ? _08097_ : _08096_;
  assign _08099_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [6] : \MSYNC_1r1w.synth.nz.mem[892] [6];
  assign _08100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [6] : \MSYNC_1r1w.synth.nz.mem[894] [6];
  assign _08101_ = \bapg_rd.w_ptr_r [1] ? _08100_ : _08099_;
  assign _08102_ = \bapg_rd.w_ptr_r [2] ? _08101_ : _08098_;
  assign _08103_ = \bapg_rd.w_ptr_r [3] ? _08102_ : _08095_;
  assign _08104_ = \bapg_rd.w_ptr_r [4] ? _08103_ : _08088_;
  assign _08105_ = \bapg_rd.w_ptr_r [5] ? _08104_ : _08073_;
  assign _08106_ = \bapg_rd.w_ptr_r [6] ? _08105_ : _08042_;
  assign _08107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [6] : \MSYNC_1r1w.synth.nz.mem[896] [6];
  assign _08108_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [6] : \MSYNC_1r1w.synth.nz.mem[898] [6];
  assign _08109_ = \bapg_rd.w_ptr_r [1] ? _08108_ : _08107_;
  assign _08110_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [6] : \MSYNC_1r1w.synth.nz.mem[900] [6];
  assign _08111_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [6] : \MSYNC_1r1w.synth.nz.mem[902] [6];
  assign _08112_ = \bapg_rd.w_ptr_r [1] ? _08111_ : _08110_;
  assign _08113_ = \bapg_rd.w_ptr_r [2] ? _08112_ : _08109_;
  assign _08114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [6] : \MSYNC_1r1w.synth.nz.mem[904] [6];
  assign _08115_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [6] : \MSYNC_1r1w.synth.nz.mem[906] [6];
  assign _08116_ = \bapg_rd.w_ptr_r [1] ? _08115_ : _08114_;
  assign _08117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [6] : \MSYNC_1r1w.synth.nz.mem[908] [6];
  assign _08118_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [6] : \MSYNC_1r1w.synth.nz.mem[910] [6];
  assign _08119_ = \bapg_rd.w_ptr_r [1] ? _08118_ : _08117_;
  assign _08120_ = \bapg_rd.w_ptr_r [2] ? _08119_ : _08116_;
  assign _08121_ = \bapg_rd.w_ptr_r [3] ? _08120_ : _08113_;
  assign _08122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [6] : \MSYNC_1r1w.synth.nz.mem[912] [6];
  assign _08123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [6] : \MSYNC_1r1w.synth.nz.mem[914] [6];
  assign _08124_ = \bapg_rd.w_ptr_r [1] ? _08123_ : _08122_;
  assign _08125_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [6] : \MSYNC_1r1w.synth.nz.mem[916] [6];
  assign _08126_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [6] : \MSYNC_1r1w.synth.nz.mem[918] [6];
  assign _08127_ = \bapg_rd.w_ptr_r [1] ? _08126_ : _08125_;
  assign _08128_ = \bapg_rd.w_ptr_r [2] ? _08127_ : _08124_;
  assign _08129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [6] : \MSYNC_1r1w.synth.nz.mem[920] [6];
  assign _08130_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [6] : \MSYNC_1r1w.synth.nz.mem[922] [6];
  assign _08131_ = \bapg_rd.w_ptr_r [1] ? _08130_ : _08129_;
  assign _08132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [6] : \MSYNC_1r1w.synth.nz.mem[924] [6];
  assign _08133_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [6] : \MSYNC_1r1w.synth.nz.mem[926] [6];
  assign _08134_ = \bapg_rd.w_ptr_r [1] ? _08133_ : _08132_;
  assign _08135_ = \bapg_rd.w_ptr_r [2] ? _08134_ : _08131_;
  assign _08136_ = \bapg_rd.w_ptr_r [3] ? _08135_ : _08128_;
  assign _08137_ = \bapg_rd.w_ptr_r [4] ? _08136_ : _08121_;
  assign _08138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [6] : \MSYNC_1r1w.synth.nz.mem[928] [6];
  assign _08139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [6] : \MSYNC_1r1w.synth.nz.mem[930] [6];
  assign _08140_ = \bapg_rd.w_ptr_r [1] ? _08139_ : _08138_;
  assign _08141_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [6] : \MSYNC_1r1w.synth.nz.mem[932] [6];
  assign _08142_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [6] : \MSYNC_1r1w.synth.nz.mem[934] [6];
  assign _08143_ = \bapg_rd.w_ptr_r [1] ? _08142_ : _08141_;
  assign _08144_ = \bapg_rd.w_ptr_r [2] ? _08143_ : _08140_;
  assign _08145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [6] : \MSYNC_1r1w.synth.nz.mem[936] [6];
  assign _08146_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [6] : \MSYNC_1r1w.synth.nz.mem[938] [6];
  assign _08147_ = \bapg_rd.w_ptr_r [1] ? _08146_ : _08145_;
  assign _08148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [6] : \MSYNC_1r1w.synth.nz.mem[940] [6];
  assign _08149_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [6] : \MSYNC_1r1w.synth.nz.mem[942] [6];
  assign _08150_ = \bapg_rd.w_ptr_r [1] ? _08149_ : _08148_;
  assign _08151_ = \bapg_rd.w_ptr_r [2] ? _08150_ : _08147_;
  assign _08152_ = \bapg_rd.w_ptr_r [3] ? _08151_ : _08144_;
  assign _08153_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [6] : \MSYNC_1r1w.synth.nz.mem[944] [6];
  assign _08154_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [6] : \MSYNC_1r1w.synth.nz.mem[946] [6];
  assign _08155_ = \bapg_rd.w_ptr_r [1] ? _08154_ : _08153_;
  assign _08156_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [6] : \MSYNC_1r1w.synth.nz.mem[948] [6];
  assign _08157_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [6] : \MSYNC_1r1w.synth.nz.mem[950] [6];
  assign _08158_ = \bapg_rd.w_ptr_r [1] ? _08157_ : _08156_;
  assign _08159_ = \bapg_rd.w_ptr_r [2] ? _08158_ : _08155_;
  assign _08160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [6] : \MSYNC_1r1w.synth.nz.mem[952] [6];
  assign _08161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [6] : \MSYNC_1r1w.synth.nz.mem[954] [6];
  assign _08162_ = \bapg_rd.w_ptr_r [1] ? _08161_ : _08160_;
  assign _08163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [6] : \MSYNC_1r1w.synth.nz.mem[956] [6];
  assign _08164_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [6] : \MSYNC_1r1w.synth.nz.mem[958] [6];
  assign _08165_ = \bapg_rd.w_ptr_r [1] ? _08164_ : _08163_;
  assign _08166_ = \bapg_rd.w_ptr_r [2] ? _08165_ : _08162_;
  assign _08167_ = \bapg_rd.w_ptr_r [3] ? _08166_ : _08159_;
  assign _08168_ = \bapg_rd.w_ptr_r [4] ? _08167_ : _08152_;
  assign _08169_ = \bapg_rd.w_ptr_r [5] ? _08168_ : _08137_;
  assign _08170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [6] : \MSYNC_1r1w.synth.nz.mem[960] [6];
  assign _08171_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [6] : \MSYNC_1r1w.synth.nz.mem[962] [6];
  assign _08172_ = \bapg_rd.w_ptr_r [1] ? _08171_ : _08170_;
  assign _08173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [6] : \MSYNC_1r1w.synth.nz.mem[964] [6];
  assign _08174_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [6] : \MSYNC_1r1w.synth.nz.mem[966] [6];
  assign _08175_ = \bapg_rd.w_ptr_r [1] ? _08174_ : _08173_;
  assign _08176_ = \bapg_rd.w_ptr_r [2] ? _08175_ : _08172_;
  assign _08177_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [6] : \MSYNC_1r1w.synth.nz.mem[968] [6];
  assign _08178_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [6] : \MSYNC_1r1w.synth.nz.mem[970] [6];
  assign _08179_ = \bapg_rd.w_ptr_r [1] ? _08178_ : _08177_;
  assign _08180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [6] : \MSYNC_1r1w.synth.nz.mem[972] [6];
  assign _08181_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [6] : \MSYNC_1r1w.synth.nz.mem[974] [6];
  assign _08182_ = \bapg_rd.w_ptr_r [1] ? _08181_ : _08180_;
  assign _08183_ = \bapg_rd.w_ptr_r [2] ? _08182_ : _08179_;
  assign _08184_ = \bapg_rd.w_ptr_r [3] ? _08183_ : _08176_;
  assign _08185_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [6] : \MSYNC_1r1w.synth.nz.mem[976] [6];
  assign _08186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [6] : \MSYNC_1r1w.synth.nz.mem[978] [6];
  assign _08187_ = \bapg_rd.w_ptr_r [1] ? _08186_ : _08185_;
  assign _08188_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [6] : \MSYNC_1r1w.synth.nz.mem[980] [6];
  assign _08189_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [6] : \MSYNC_1r1w.synth.nz.mem[982] [6];
  assign _08190_ = \bapg_rd.w_ptr_r [1] ? _08189_ : _08188_;
  assign _08191_ = \bapg_rd.w_ptr_r [2] ? _08190_ : _08187_;
  assign _08192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [6] : \MSYNC_1r1w.synth.nz.mem[984] [6];
  assign _08193_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [6] : \MSYNC_1r1w.synth.nz.mem[986] [6];
  assign _08194_ = \bapg_rd.w_ptr_r [1] ? _08193_ : _08192_;
  assign _08195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [6] : \MSYNC_1r1w.synth.nz.mem[988] [6];
  assign _08196_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [6] : \MSYNC_1r1w.synth.nz.mem[990] [6];
  assign _08197_ = \bapg_rd.w_ptr_r [1] ? _08196_ : _08195_;
  assign _08198_ = \bapg_rd.w_ptr_r [2] ? _08197_ : _08194_;
  assign _08199_ = \bapg_rd.w_ptr_r [3] ? _08198_ : _08191_;
  assign _08200_ = \bapg_rd.w_ptr_r [4] ? _08199_ : _08184_;
  assign _08201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [6] : \MSYNC_1r1w.synth.nz.mem[992] [6];
  assign _08202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [6] : \MSYNC_1r1w.synth.nz.mem[994] [6];
  assign _08203_ = \bapg_rd.w_ptr_r [1] ? _08202_ : _08201_;
  assign _08204_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [6] : \MSYNC_1r1w.synth.nz.mem[996] [6];
  assign _08205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [6] : \MSYNC_1r1w.synth.nz.mem[998] [6];
  assign _08206_ = \bapg_rd.w_ptr_r [1] ? _08205_ : _08204_;
  assign _08207_ = \bapg_rd.w_ptr_r [2] ? _08206_ : _08203_;
  assign _08208_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [6] : \MSYNC_1r1w.synth.nz.mem[1000] [6];
  assign _08209_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [6] : \MSYNC_1r1w.synth.nz.mem[1002] [6];
  assign _08210_ = \bapg_rd.w_ptr_r [1] ? _08209_ : _08208_;
  assign _08211_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [6] : \MSYNC_1r1w.synth.nz.mem[1004] [6];
  assign _08212_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [6] : \MSYNC_1r1w.synth.nz.mem[1006] [6];
  assign _08213_ = \bapg_rd.w_ptr_r [1] ? _08212_ : _08211_;
  assign _08214_ = \bapg_rd.w_ptr_r [2] ? _08213_ : _08210_;
  assign _08215_ = \bapg_rd.w_ptr_r [3] ? _08214_ : _08207_;
  assign _08216_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [6] : \MSYNC_1r1w.synth.nz.mem[1008] [6];
  assign _08217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [6] : \MSYNC_1r1w.synth.nz.mem[1010] [6];
  assign _08218_ = \bapg_rd.w_ptr_r [1] ? _08217_ : _08216_;
  assign _08219_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [6] : \MSYNC_1r1w.synth.nz.mem[1012] [6];
  assign _08220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [6] : \MSYNC_1r1w.synth.nz.mem[1014] [6];
  assign _08221_ = \bapg_rd.w_ptr_r [1] ? _08220_ : _08219_;
  assign _08222_ = \bapg_rd.w_ptr_r [2] ? _08221_ : _08218_;
  assign _08223_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [6] : \MSYNC_1r1w.synth.nz.mem[1016] [6];
  assign _08224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [6] : \MSYNC_1r1w.synth.nz.mem[1018] [6];
  assign _08225_ = \bapg_rd.w_ptr_r [1] ? _08224_ : _08223_;
  assign _08226_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [6] : \MSYNC_1r1w.synth.nz.mem[1020] [6];
  assign _08227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [6] : \MSYNC_1r1w.synth.nz.mem[1022] [6];
  assign _08228_ = \bapg_rd.w_ptr_r [1] ? _08227_ : _08226_;
  assign _08229_ = \bapg_rd.w_ptr_r [2] ? _08228_ : _08225_;
  assign _08230_ = \bapg_rd.w_ptr_r [3] ? _08229_ : _08222_;
  assign _08231_ = \bapg_rd.w_ptr_r [4] ? _08230_ : _08215_;
  assign _08232_ = \bapg_rd.w_ptr_r [5] ? _08231_ : _08200_;
  assign _08233_ = \bapg_rd.w_ptr_r [6] ? _08232_ : _08169_;
  assign _08234_ = \bapg_rd.w_ptr_r [7] ? _08233_ : _08106_;
  assign _08235_ = \bapg_rd.w_ptr_r [8] ? _08234_ : _07979_;
  assign r_data_o[6] = \bapg_rd.w_ptr_r [9] ? _08235_ : _07724_;
  assign _08236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [7] : \MSYNC_1r1w.synth.nz.mem[0] [7];
  assign _08237_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [7] : \MSYNC_1r1w.synth.nz.mem[2] [7];
  assign _08238_ = \bapg_rd.w_ptr_r [1] ? _08237_ : _08236_;
  assign _08239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [7] : \MSYNC_1r1w.synth.nz.mem[4] [7];
  assign _08240_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [7] : \MSYNC_1r1w.synth.nz.mem[6] [7];
  assign _08241_ = \bapg_rd.w_ptr_r [1] ? _08240_ : _08239_;
  assign _08242_ = \bapg_rd.w_ptr_r [2] ? _08241_ : _08238_;
  assign _08243_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [7] : \MSYNC_1r1w.synth.nz.mem[8] [7];
  assign _08244_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [7] : \MSYNC_1r1w.synth.nz.mem[10] [7];
  assign _08245_ = \bapg_rd.w_ptr_r [1] ? _08244_ : _08243_;
  assign _08246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [7] : \MSYNC_1r1w.synth.nz.mem[12] [7];
  assign _08247_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [7] : \MSYNC_1r1w.synth.nz.mem[14] [7];
  assign _08248_ = \bapg_rd.w_ptr_r [1] ? _08247_ : _08246_;
  assign _08249_ = \bapg_rd.w_ptr_r [2] ? _08248_ : _08245_;
  assign _08250_ = \bapg_rd.w_ptr_r [3] ? _08249_ : _08242_;
  assign _08251_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [7] : \MSYNC_1r1w.synth.nz.mem[16] [7];
  assign _08252_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [7] : \MSYNC_1r1w.synth.nz.mem[18] [7];
  assign _08253_ = \bapg_rd.w_ptr_r [1] ? _08252_ : _08251_;
  assign _08254_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [7] : \MSYNC_1r1w.synth.nz.mem[20] [7];
  assign _08255_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [7] : \MSYNC_1r1w.synth.nz.mem[22] [7];
  assign _08256_ = \bapg_rd.w_ptr_r [1] ? _08255_ : _08254_;
  assign _08257_ = \bapg_rd.w_ptr_r [2] ? _08256_ : _08253_;
  assign _08258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [7] : \MSYNC_1r1w.synth.nz.mem[24] [7];
  assign _08259_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [7] : \MSYNC_1r1w.synth.nz.mem[26] [7];
  assign _08260_ = \bapg_rd.w_ptr_r [1] ? _08259_ : _08258_;
  assign _08261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [7] : \MSYNC_1r1w.synth.nz.mem[28] [7];
  assign _08262_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [7] : \MSYNC_1r1w.synth.nz.mem[30] [7];
  assign _08263_ = \bapg_rd.w_ptr_r [1] ? _08262_ : _08261_;
  assign _08264_ = \bapg_rd.w_ptr_r [2] ? _08263_ : _08260_;
  assign _08265_ = \bapg_rd.w_ptr_r [3] ? _08264_ : _08257_;
  assign _08266_ = \bapg_rd.w_ptr_r [4] ? _08265_ : _08250_;
  assign _08267_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [7] : \MSYNC_1r1w.synth.nz.mem[32] [7];
  assign _08268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [7] : \MSYNC_1r1w.synth.nz.mem[34] [7];
  assign _08269_ = \bapg_rd.w_ptr_r [1] ? _08268_ : _08267_;
  assign _08270_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [7] : \MSYNC_1r1w.synth.nz.mem[36] [7];
  assign _08271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [7] : \MSYNC_1r1w.synth.nz.mem[38] [7];
  assign _08272_ = \bapg_rd.w_ptr_r [1] ? _08271_ : _08270_;
  assign _08273_ = \bapg_rd.w_ptr_r [2] ? _08272_ : _08269_;
  assign _08274_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [7] : \MSYNC_1r1w.synth.nz.mem[40] [7];
  assign _08275_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [7] : \MSYNC_1r1w.synth.nz.mem[42] [7];
  assign _08276_ = \bapg_rd.w_ptr_r [1] ? _08275_ : _08274_;
  assign _08277_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [7] : \MSYNC_1r1w.synth.nz.mem[44] [7];
  assign _08278_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [7] : \MSYNC_1r1w.synth.nz.mem[46] [7];
  assign _08279_ = \bapg_rd.w_ptr_r [1] ? _08278_ : _08277_;
  assign _08280_ = \bapg_rd.w_ptr_r [2] ? _08279_ : _08276_;
  assign _08281_ = \bapg_rd.w_ptr_r [3] ? _08280_ : _08273_;
  assign _08282_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [7] : \MSYNC_1r1w.synth.nz.mem[48] [7];
  assign _08283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [7] : \MSYNC_1r1w.synth.nz.mem[50] [7];
  assign _08284_ = \bapg_rd.w_ptr_r [1] ? _08283_ : _08282_;
  assign _08285_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [7] : \MSYNC_1r1w.synth.nz.mem[52] [7];
  assign _08286_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [7] : \MSYNC_1r1w.synth.nz.mem[54] [7];
  assign _08287_ = \bapg_rd.w_ptr_r [1] ? _08286_ : _08285_;
  assign _08288_ = \bapg_rd.w_ptr_r [2] ? _08287_ : _08284_;
  assign _08289_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [7] : \MSYNC_1r1w.synth.nz.mem[56] [7];
  assign _08290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [7] : \MSYNC_1r1w.synth.nz.mem[58] [7];
  assign _08291_ = \bapg_rd.w_ptr_r [1] ? _08290_ : _08289_;
  assign _08292_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [7] : \MSYNC_1r1w.synth.nz.mem[60] [7];
  assign _08293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [7] : \MSYNC_1r1w.synth.nz.mem[62] [7];
  assign _08294_ = \bapg_rd.w_ptr_r [1] ? _08293_ : _08292_;
  assign _08295_ = \bapg_rd.w_ptr_r [2] ? _08294_ : _08291_;
  assign _08296_ = \bapg_rd.w_ptr_r [3] ? _08295_ : _08288_;
  assign _08297_ = \bapg_rd.w_ptr_r [4] ? _08296_ : _08281_;
  assign _08298_ = \bapg_rd.w_ptr_r [5] ? _08297_ : _08266_;
  assign _08299_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [7] : \MSYNC_1r1w.synth.nz.mem[64] [7];
  assign _08300_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [7] : \MSYNC_1r1w.synth.nz.mem[66] [7];
  assign _08301_ = \bapg_rd.w_ptr_r [1] ? _08300_ : _08299_;
  assign _08302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [7] : \MSYNC_1r1w.synth.nz.mem[68] [7];
  assign _08303_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [7] : \MSYNC_1r1w.synth.nz.mem[70] [7];
  assign _08304_ = \bapg_rd.w_ptr_r [1] ? _08303_ : _08302_;
  assign _08305_ = \bapg_rd.w_ptr_r [2] ? _08304_ : _08301_;
  assign _08306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [7] : \MSYNC_1r1w.synth.nz.mem[72] [7];
  assign _08307_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [7] : \MSYNC_1r1w.synth.nz.mem[74] [7];
  assign _08308_ = \bapg_rd.w_ptr_r [1] ? _08307_ : _08306_;
  assign _08309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [7] : \MSYNC_1r1w.synth.nz.mem[76] [7];
  assign _08310_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [7] : \MSYNC_1r1w.synth.nz.mem[78] [7];
  assign _08311_ = \bapg_rd.w_ptr_r [1] ? _08310_ : _08309_;
  assign _08312_ = \bapg_rd.w_ptr_r [2] ? _08311_ : _08308_;
  assign _08313_ = \bapg_rd.w_ptr_r [3] ? _08312_ : _08305_;
  assign _08314_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [7] : \MSYNC_1r1w.synth.nz.mem[80] [7];
  assign _08315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [7] : \MSYNC_1r1w.synth.nz.mem[82] [7];
  assign _08316_ = \bapg_rd.w_ptr_r [1] ? _08315_ : _08314_;
  assign _08317_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [7] : \MSYNC_1r1w.synth.nz.mem[84] [7];
  assign _08318_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [7] : \MSYNC_1r1w.synth.nz.mem[86] [7];
  assign _08319_ = \bapg_rd.w_ptr_r [1] ? _08318_ : _08317_;
  assign _08320_ = \bapg_rd.w_ptr_r [2] ? _08319_ : _08316_;
  assign _08321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [7] : \MSYNC_1r1w.synth.nz.mem[88] [7];
  assign _08322_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [7] : \MSYNC_1r1w.synth.nz.mem[90] [7];
  assign _08323_ = \bapg_rd.w_ptr_r [1] ? _08322_ : _08321_;
  assign _08324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [7] : \MSYNC_1r1w.synth.nz.mem[92] [7];
  assign _08325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [7] : \MSYNC_1r1w.synth.nz.mem[94] [7];
  assign _08326_ = \bapg_rd.w_ptr_r [1] ? _08325_ : _08324_;
  assign _08327_ = \bapg_rd.w_ptr_r [2] ? _08326_ : _08323_;
  assign _08328_ = \bapg_rd.w_ptr_r [3] ? _08327_ : _08320_;
  assign _08329_ = \bapg_rd.w_ptr_r [4] ? _08328_ : _08313_;
  assign _08330_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [7] : \MSYNC_1r1w.synth.nz.mem[96] [7];
  assign _08331_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [7] : \MSYNC_1r1w.synth.nz.mem[98] [7];
  assign _08332_ = \bapg_rd.w_ptr_r [1] ? _08331_ : _08330_;
  assign _08333_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [7] : \MSYNC_1r1w.synth.nz.mem[100] [7];
  assign _08334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [7] : \MSYNC_1r1w.synth.nz.mem[102] [7];
  assign _08335_ = \bapg_rd.w_ptr_r [1] ? _08334_ : _08333_;
  assign _08336_ = \bapg_rd.w_ptr_r [2] ? _08335_ : _08332_;
  assign _08337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [7] : \MSYNC_1r1w.synth.nz.mem[104] [7];
  assign _08338_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [7] : \MSYNC_1r1w.synth.nz.mem[106] [7];
  assign _08339_ = \bapg_rd.w_ptr_r [1] ? _08338_ : _08337_;
  assign _08340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [7] : \MSYNC_1r1w.synth.nz.mem[108] [7];
  assign _08341_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [7] : \MSYNC_1r1w.synth.nz.mem[110] [7];
  assign _08342_ = \bapg_rd.w_ptr_r [1] ? _08341_ : _08340_;
  assign _08343_ = \bapg_rd.w_ptr_r [2] ? _08342_ : _08339_;
  assign _08344_ = \bapg_rd.w_ptr_r [3] ? _08343_ : _08336_;
  assign _08345_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [7] : \MSYNC_1r1w.synth.nz.mem[112] [7];
  assign _08346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [7] : \MSYNC_1r1w.synth.nz.mem[114] [7];
  assign _08347_ = \bapg_rd.w_ptr_r [1] ? _08346_ : _08345_;
  assign _08348_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [7] : \MSYNC_1r1w.synth.nz.mem[116] [7];
  assign _08349_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [7] : \MSYNC_1r1w.synth.nz.mem[118] [7];
  assign _08350_ = \bapg_rd.w_ptr_r [1] ? _08349_ : _08348_;
  assign _08351_ = \bapg_rd.w_ptr_r [2] ? _08350_ : _08347_;
  assign _08352_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [7] : \MSYNC_1r1w.synth.nz.mem[120] [7];
  assign _08353_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [7] : \MSYNC_1r1w.synth.nz.mem[122] [7];
  assign _08354_ = \bapg_rd.w_ptr_r [1] ? _08353_ : _08352_;
  assign _08355_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [7] : \MSYNC_1r1w.synth.nz.mem[124] [7];
  assign _08356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [7] : \MSYNC_1r1w.synth.nz.mem[126] [7];
  assign _08357_ = \bapg_rd.w_ptr_r [1] ? _08356_ : _08355_;
  assign _08358_ = \bapg_rd.w_ptr_r [2] ? _08357_ : _08354_;
  assign _08359_ = \bapg_rd.w_ptr_r [3] ? _08358_ : _08351_;
  assign _08360_ = \bapg_rd.w_ptr_r [4] ? _08359_ : _08344_;
  assign _08361_ = \bapg_rd.w_ptr_r [5] ? _08360_ : _08329_;
  assign _08362_ = \bapg_rd.w_ptr_r [6] ? _08361_ : _08298_;
  assign _08363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [7] : \MSYNC_1r1w.synth.nz.mem[128] [7];
  assign _08364_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [7] : \MSYNC_1r1w.synth.nz.mem[130] [7];
  assign _08365_ = \bapg_rd.w_ptr_r [1] ? _08364_ : _08363_;
  assign _08366_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [7] : \MSYNC_1r1w.synth.nz.mem[132] [7];
  assign _08367_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [7] : \MSYNC_1r1w.synth.nz.mem[134] [7];
  assign _08368_ = \bapg_rd.w_ptr_r [1] ? _08367_ : _08366_;
  assign _08369_ = \bapg_rd.w_ptr_r [2] ? _08368_ : _08365_;
  assign _08370_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [7] : \MSYNC_1r1w.synth.nz.mem[136] [7];
  assign _08371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [7] : \MSYNC_1r1w.synth.nz.mem[138] [7];
  assign _08372_ = \bapg_rd.w_ptr_r [1] ? _08371_ : _08370_;
  assign _08373_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [7] : \MSYNC_1r1w.synth.nz.mem[140] [7];
  assign _08374_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [7] : \MSYNC_1r1w.synth.nz.mem[142] [7];
  assign _08375_ = \bapg_rd.w_ptr_r [1] ? _08374_ : _08373_;
  assign _08376_ = \bapg_rd.w_ptr_r [2] ? _08375_ : _08372_;
  assign _08377_ = \bapg_rd.w_ptr_r [3] ? _08376_ : _08369_;
  assign _08378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [7] : \MSYNC_1r1w.synth.nz.mem[144] [7];
  assign _08379_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [7] : \MSYNC_1r1w.synth.nz.mem[146] [7];
  assign _08380_ = \bapg_rd.w_ptr_r [1] ? _08379_ : _08378_;
  assign _08381_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [7] : \MSYNC_1r1w.synth.nz.mem[148] [7];
  assign _08382_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [7] : \MSYNC_1r1w.synth.nz.mem[150] [7];
  assign _08383_ = \bapg_rd.w_ptr_r [1] ? _08382_ : _08381_;
  assign _08384_ = \bapg_rd.w_ptr_r [2] ? _08383_ : _08380_;
  assign _08385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [7] : \MSYNC_1r1w.synth.nz.mem[152] [7];
  assign _08386_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [7] : \MSYNC_1r1w.synth.nz.mem[154] [7];
  assign _08387_ = \bapg_rd.w_ptr_r [1] ? _08386_ : _08385_;
  assign _08388_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [7] : \MSYNC_1r1w.synth.nz.mem[156] [7];
  assign _08389_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [7] : \MSYNC_1r1w.synth.nz.mem[158] [7];
  assign _08390_ = \bapg_rd.w_ptr_r [1] ? _08389_ : _08388_;
  assign _08391_ = \bapg_rd.w_ptr_r [2] ? _08390_ : _08387_;
  assign _08392_ = \bapg_rd.w_ptr_r [3] ? _08391_ : _08384_;
  assign _08393_ = \bapg_rd.w_ptr_r [4] ? _08392_ : _08377_;
  assign _08394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [7] : \MSYNC_1r1w.synth.nz.mem[160] [7];
  assign _08395_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [7] : \MSYNC_1r1w.synth.nz.mem[162] [7];
  assign _08396_ = \bapg_rd.w_ptr_r [1] ? _08395_ : _08394_;
  assign _08397_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [7] : \MSYNC_1r1w.synth.nz.mem[164] [7];
  assign _08398_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [7] : \MSYNC_1r1w.synth.nz.mem[166] [7];
  assign _08399_ = \bapg_rd.w_ptr_r [1] ? _08398_ : _08397_;
  assign _08400_ = \bapg_rd.w_ptr_r [2] ? _08399_ : _08396_;
  assign _08401_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [7] : \MSYNC_1r1w.synth.nz.mem[168] [7];
  assign _08402_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [7] : \MSYNC_1r1w.synth.nz.mem[170] [7];
  assign _08403_ = \bapg_rd.w_ptr_r [1] ? _08402_ : _08401_;
  assign _08404_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [7] : \MSYNC_1r1w.synth.nz.mem[172] [7];
  assign _08405_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [7] : \MSYNC_1r1w.synth.nz.mem[174] [7];
  assign _08406_ = \bapg_rd.w_ptr_r [1] ? _08405_ : _08404_;
  assign _08407_ = \bapg_rd.w_ptr_r [2] ? _08406_ : _08403_;
  assign _08408_ = \bapg_rd.w_ptr_r [3] ? _08407_ : _08400_;
  assign _08409_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [7] : \MSYNC_1r1w.synth.nz.mem[176] [7];
  assign _08410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [7] : \MSYNC_1r1w.synth.nz.mem[178] [7];
  assign _08411_ = \bapg_rd.w_ptr_r [1] ? _08410_ : _08409_;
  assign _08412_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [7] : \MSYNC_1r1w.synth.nz.mem[180] [7];
  assign _08413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [7] : \MSYNC_1r1w.synth.nz.mem[182] [7];
  assign _08414_ = \bapg_rd.w_ptr_r [1] ? _08413_ : _08412_;
  assign _08415_ = \bapg_rd.w_ptr_r [2] ? _08414_ : _08411_;
  assign _08416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [7] : \MSYNC_1r1w.synth.nz.mem[184] [7];
  assign _08417_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [7] : \MSYNC_1r1w.synth.nz.mem[186] [7];
  assign _08418_ = \bapg_rd.w_ptr_r [1] ? _08417_ : _08416_;
  assign _08419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [7] : \MSYNC_1r1w.synth.nz.mem[188] [7];
  assign _08420_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [7] : \MSYNC_1r1w.synth.nz.mem[190] [7];
  assign _08421_ = \bapg_rd.w_ptr_r [1] ? _08420_ : _08419_;
  assign _08422_ = \bapg_rd.w_ptr_r [2] ? _08421_ : _08418_;
  assign _08423_ = \bapg_rd.w_ptr_r [3] ? _08422_ : _08415_;
  assign _08424_ = \bapg_rd.w_ptr_r [4] ? _08423_ : _08408_;
  assign _08425_ = \bapg_rd.w_ptr_r [5] ? _08424_ : _08393_;
  assign _08426_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [7] : \MSYNC_1r1w.synth.nz.mem[192] [7];
  assign _08427_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [7] : \MSYNC_1r1w.synth.nz.mem[194] [7];
  assign _08428_ = \bapg_rd.w_ptr_r [1] ? _08427_ : _08426_;
  assign _08429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [7] : \MSYNC_1r1w.synth.nz.mem[196] [7];
  assign _08430_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [7] : \MSYNC_1r1w.synth.nz.mem[198] [7];
  assign _08431_ = \bapg_rd.w_ptr_r [1] ? _08430_ : _08429_;
  assign _08432_ = \bapg_rd.w_ptr_r [2] ? _08431_ : _08428_;
  assign _08433_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [7] : \MSYNC_1r1w.synth.nz.mem[200] [7];
  assign _08434_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [7] : \MSYNC_1r1w.synth.nz.mem[202] [7];
  assign _08435_ = \bapg_rd.w_ptr_r [1] ? _08434_ : _08433_;
  assign _08436_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [7] : \MSYNC_1r1w.synth.nz.mem[204] [7];
  assign _08437_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [7] : \MSYNC_1r1w.synth.nz.mem[206] [7];
  assign _08438_ = \bapg_rd.w_ptr_r [1] ? _08437_ : _08436_;
  assign _08439_ = \bapg_rd.w_ptr_r [2] ? _08438_ : _08435_;
  assign _08440_ = \bapg_rd.w_ptr_r [3] ? _08439_ : _08432_;
  assign _08441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [7] : \MSYNC_1r1w.synth.nz.mem[208] [7];
  assign _08442_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [7] : \MSYNC_1r1w.synth.nz.mem[210] [7];
  assign _08443_ = \bapg_rd.w_ptr_r [1] ? _08442_ : _08441_;
  assign _08444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [7] : \MSYNC_1r1w.synth.nz.mem[212] [7];
  assign _08445_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [7] : \MSYNC_1r1w.synth.nz.mem[214] [7];
  assign _08446_ = \bapg_rd.w_ptr_r [1] ? _08445_ : _08444_;
  assign _08447_ = \bapg_rd.w_ptr_r [2] ? _08446_ : _08443_;
  assign _08448_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [7] : \MSYNC_1r1w.synth.nz.mem[216] [7];
  assign _08449_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [7] : \MSYNC_1r1w.synth.nz.mem[218] [7];
  assign _08450_ = \bapg_rd.w_ptr_r [1] ? _08449_ : _08448_;
  assign _08451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [7] : \MSYNC_1r1w.synth.nz.mem[220] [7];
  assign _08452_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [7] : \MSYNC_1r1w.synth.nz.mem[222] [7];
  assign _08453_ = \bapg_rd.w_ptr_r [1] ? _08452_ : _08451_;
  assign _08454_ = \bapg_rd.w_ptr_r [2] ? _08453_ : _08450_;
  assign _08455_ = \bapg_rd.w_ptr_r [3] ? _08454_ : _08447_;
  assign _08456_ = \bapg_rd.w_ptr_r [4] ? _08455_ : _08440_;
  assign _08457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [7] : \MSYNC_1r1w.synth.nz.mem[224] [7];
  assign _08458_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [7] : \MSYNC_1r1w.synth.nz.mem[226] [7];
  assign _08459_ = \bapg_rd.w_ptr_r [1] ? _08458_ : _08457_;
  assign _08460_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [7] : \MSYNC_1r1w.synth.nz.mem[228] [7];
  assign _08461_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [7] : \MSYNC_1r1w.synth.nz.mem[230] [7];
  assign _08462_ = \bapg_rd.w_ptr_r [1] ? _08461_ : _08460_;
  assign _08463_ = \bapg_rd.w_ptr_r [2] ? _08462_ : _08459_;
  assign _08464_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [7] : \MSYNC_1r1w.synth.nz.mem[232] [7];
  assign _08465_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [7] : \MSYNC_1r1w.synth.nz.mem[234] [7];
  assign _08466_ = \bapg_rd.w_ptr_r [1] ? _08465_ : _08464_;
  assign _08467_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [7] : \MSYNC_1r1w.synth.nz.mem[236] [7];
  assign _08468_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [7] : \MSYNC_1r1w.synth.nz.mem[238] [7];
  assign _08469_ = \bapg_rd.w_ptr_r [1] ? _08468_ : _08467_;
  assign _08470_ = \bapg_rd.w_ptr_r [2] ? _08469_ : _08466_;
  assign _08471_ = \bapg_rd.w_ptr_r [3] ? _08470_ : _08463_;
  assign _08472_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [7] : \MSYNC_1r1w.synth.nz.mem[240] [7];
  assign _08473_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [7] : \MSYNC_1r1w.synth.nz.mem[242] [7];
  assign _08474_ = \bapg_rd.w_ptr_r [1] ? _08473_ : _08472_;
  assign _08475_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [7] : \MSYNC_1r1w.synth.nz.mem[244] [7];
  assign _08476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [7] : \MSYNC_1r1w.synth.nz.mem[246] [7];
  assign _08477_ = \bapg_rd.w_ptr_r [1] ? _08476_ : _08475_;
  assign _08478_ = \bapg_rd.w_ptr_r [2] ? _08477_ : _08474_;
  assign _08479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [7] : \MSYNC_1r1w.synth.nz.mem[248] [7];
  assign _08480_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [7] : \MSYNC_1r1w.synth.nz.mem[250] [7];
  assign _08481_ = \bapg_rd.w_ptr_r [1] ? _08480_ : _08479_;
  assign _08482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [7] : \MSYNC_1r1w.synth.nz.mem[252] [7];
  assign _08483_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [7] : \MSYNC_1r1w.synth.nz.mem[254] [7];
  assign _08484_ = \bapg_rd.w_ptr_r [1] ? _08483_ : _08482_;
  assign _08485_ = \bapg_rd.w_ptr_r [2] ? _08484_ : _08481_;
  assign _08486_ = \bapg_rd.w_ptr_r [3] ? _08485_ : _08478_;
  assign _08487_ = \bapg_rd.w_ptr_r [4] ? _08486_ : _08471_;
  assign _08488_ = \bapg_rd.w_ptr_r [5] ? _08487_ : _08456_;
  assign _08489_ = \bapg_rd.w_ptr_r [6] ? _08488_ : _08425_;
  assign _08490_ = \bapg_rd.w_ptr_r [7] ? _08489_ : _08362_;
  assign _08491_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [7] : \MSYNC_1r1w.synth.nz.mem[256] [7];
  assign _08492_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [7] : \MSYNC_1r1w.synth.nz.mem[258] [7];
  assign _08493_ = \bapg_rd.w_ptr_r [1] ? _08492_ : _08491_;
  assign _08494_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [7] : \MSYNC_1r1w.synth.nz.mem[260] [7];
  assign _08495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [7] : \MSYNC_1r1w.synth.nz.mem[262] [7];
  assign _08496_ = \bapg_rd.w_ptr_r [1] ? _08495_ : _08494_;
  assign _08497_ = \bapg_rd.w_ptr_r [2] ? _08496_ : _08493_;
  assign _08498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [7] : \MSYNC_1r1w.synth.nz.mem[264] [7];
  assign _08499_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [7] : \MSYNC_1r1w.synth.nz.mem[266] [7];
  assign _08500_ = \bapg_rd.w_ptr_r [1] ? _08499_ : _08498_;
  assign _08501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [7] : \MSYNC_1r1w.synth.nz.mem[268] [7];
  assign _08502_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [7] : \MSYNC_1r1w.synth.nz.mem[270] [7];
  assign _08503_ = \bapg_rd.w_ptr_r [1] ? _08502_ : _08501_;
  assign _08504_ = \bapg_rd.w_ptr_r [2] ? _08503_ : _08500_;
  assign _08505_ = \bapg_rd.w_ptr_r [3] ? _08504_ : _08497_;
  assign _08506_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [7] : \MSYNC_1r1w.synth.nz.mem[272] [7];
  assign _08507_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [7] : \MSYNC_1r1w.synth.nz.mem[274] [7];
  assign _08508_ = \bapg_rd.w_ptr_r [1] ? _08507_ : _08506_;
  assign _08509_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [7] : \MSYNC_1r1w.synth.nz.mem[276] [7];
  assign _08510_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [7] : \MSYNC_1r1w.synth.nz.mem[278] [7];
  assign _08511_ = \bapg_rd.w_ptr_r [1] ? _08510_ : _08509_;
  assign _08512_ = \bapg_rd.w_ptr_r [2] ? _08511_ : _08508_;
  assign _08513_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [7] : \MSYNC_1r1w.synth.nz.mem[280] [7];
  assign _08514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [7] : \MSYNC_1r1w.synth.nz.mem[282] [7];
  assign _08515_ = \bapg_rd.w_ptr_r [1] ? _08514_ : _08513_;
  assign _08516_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [7] : \MSYNC_1r1w.synth.nz.mem[284] [7];
  assign _08517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [7] : \MSYNC_1r1w.synth.nz.mem[286] [7];
  assign _08518_ = \bapg_rd.w_ptr_r [1] ? _08517_ : _08516_;
  assign _08519_ = \bapg_rd.w_ptr_r [2] ? _08518_ : _08515_;
  assign _08520_ = \bapg_rd.w_ptr_r [3] ? _08519_ : _08512_;
  assign _08521_ = \bapg_rd.w_ptr_r [4] ? _08520_ : _08505_;
  assign _08522_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [7] : \MSYNC_1r1w.synth.nz.mem[288] [7];
  assign _08523_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [7] : \MSYNC_1r1w.synth.nz.mem[290] [7];
  assign _08524_ = \bapg_rd.w_ptr_r [1] ? _08523_ : _08522_;
  assign _08525_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [7] : \MSYNC_1r1w.synth.nz.mem[292] [7];
  assign _08526_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [7] : \MSYNC_1r1w.synth.nz.mem[294] [7];
  assign _08527_ = \bapg_rd.w_ptr_r [1] ? _08526_ : _08525_;
  assign _08528_ = \bapg_rd.w_ptr_r [2] ? _08527_ : _08524_;
  assign _08529_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [7] : \MSYNC_1r1w.synth.nz.mem[296] [7];
  assign _08530_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [7] : \MSYNC_1r1w.synth.nz.mem[298] [7];
  assign _08531_ = \bapg_rd.w_ptr_r [1] ? _08530_ : _08529_;
  assign _08532_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [7] : \MSYNC_1r1w.synth.nz.mem[300] [7];
  assign _08533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [7] : \MSYNC_1r1w.synth.nz.mem[302] [7];
  assign _08534_ = \bapg_rd.w_ptr_r [1] ? _08533_ : _08532_;
  assign _08535_ = \bapg_rd.w_ptr_r [2] ? _08534_ : _08531_;
  assign _08536_ = \bapg_rd.w_ptr_r [3] ? _08535_ : _08528_;
  assign _08537_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [7] : \MSYNC_1r1w.synth.nz.mem[304] [7];
  assign _08538_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [7] : \MSYNC_1r1w.synth.nz.mem[306] [7];
  assign _08539_ = \bapg_rd.w_ptr_r [1] ? _08538_ : _08537_;
  assign _08540_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [7] : \MSYNC_1r1w.synth.nz.mem[308] [7];
  assign _08541_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [7] : \MSYNC_1r1w.synth.nz.mem[310] [7];
  assign _08542_ = \bapg_rd.w_ptr_r [1] ? _08541_ : _08540_;
  assign _08543_ = \bapg_rd.w_ptr_r [2] ? _08542_ : _08539_;
  assign _08544_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [7] : \MSYNC_1r1w.synth.nz.mem[312] [7];
  assign _08545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [7] : \MSYNC_1r1w.synth.nz.mem[314] [7];
  assign _08546_ = \bapg_rd.w_ptr_r [1] ? _08545_ : _08544_;
  assign _08547_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [7] : \MSYNC_1r1w.synth.nz.mem[316] [7];
  assign _08548_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [7] : \MSYNC_1r1w.synth.nz.mem[318] [7];
  assign _08549_ = \bapg_rd.w_ptr_r [1] ? _08548_ : _08547_;
  assign _08550_ = \bapg_rd.w_ptr_r [2] ? _08549_ : _08546_;
  assign _08551_ = \bapg_rd.w_ptr_r [3] ? _08550_ : _08543_;
  assign _08552_ = \bapg_rd.w_ptr_r [4] ? _08551_ : _08536_;
  assign _08553_ = \bapg_rd.w_ptr_r [5] ? _08552_ : _08521_;
  assign _08554_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [7] : \MSYNC_1r1w.synth.nz.mem[320] [7];
  assign _08555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [7] : \MSYNC_1r1w.synth.nz.mem[322] [7];
  assign _08556_ = \bapg_rd.w_ptr_r [1] ? _08555_ : _08554_;
  assign _08557_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [7] : \MSYNC_1r1w.synth.nz.mem[324] [7];
  assign _08558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [7] : \MSYNC_1r1w.synth.nz.mem[326] [7];
  assign _08559_ = \bapg_rd.w_ptr_r [1] ? _08558_ : _08557_;
  assign _08560_ = \bapg_rd.w_ptr_r [2] ? _08559_ : _08556_;
  assign _08561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [7] : \MSYNC_1r1w.synth.nz.mem[328] [7];
  assign _08562_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [7] : \MSYNC_1r1w.synth.nz.mem[330] [7];
  assign _08563_ = \bapg_rd.w_ptr_r [1] ? _08562_ : _08561_;
  assign _08564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [7] : \MSYNC_1r1w.synth.nz.mem[332] [7];
  assign _08565_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [7] : \MSYNC_1r1w.synth.nz.mem[334] [7];
  assign _08566_ = \bapg_rd.w_ptr_r [1] ? _08565_ : _08564_;
  assign _08567_ = \bapg_rd.w_ptr_r [2] ? _08566_ : _08563_;
  assign _08568_ = \bapg_rd.w_ptr_r [3] ? _08567_ : _08560_;
  assign _08569_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [7] : \MSYNC_1r1w.synth.nz.mem[336] [7];
  assign _08570_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [7] : \MSYNC_1r1w.synth.nz.mem[338] [7];
  assign _08571_ = \bapg_rd.w_ptr_r [1] ? _08570_ : _08569_;
  assign _08572_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [7] : \MSYNC_1r1w.synth.nz.mem[340] [7];
  assign _08573_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [7] : \MSYNC_1r1w.synth.nz.mem[342] [7];
  assign _08574_ = \bapg_rd.w_ptr_r [1] ? _08573_ : _08572_;
  assign _08575_ = \bapg_rd.w_ptr_r [2] ? _08574_ : _08571_;
  assign _08576_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [7] : \MSYNC_1r1w.synth.nz.mem[344] [7];
  assign _08577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [7] : \MSYNC_1r1w.synth.nz.mem[346] [7];
  assign _08578_ = \bapg_rd.w_ptr_r [1] ? _08577_ : _08576_;
  assign _08579_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [7] : \MSYNC_1r1w.synth.nz.mem[348] [7];
  assign _08580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [7] : \MSYNC_1r1w.synth.nz.mem[350] [7];
  assign _08581_ = \bapg_rd.w_ptr_r [1] ? _08580_ : _08579_;
  assign _08582_ = \bapg_rd.w_ptr_r [2] ? _08581_ : _08578_;
  assign _08583_ = \bapg_rd.w_ptr_r [3] ? _08582_ : _08575_;
  assign _08584_ = \bapg_rd.w_ptr_r [4] ? _08583_ : _08568_;
  assign _08585_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [7] : \MSYNC_1r1w.synth.nz.mem[352] [7];
  assign _08586_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [7] : \MSYNC_1r1w.synth.nz.mem[354] [7];
  assign _08587_ = \bapg_rd.w_ptr_r [1] ? _08586_ : _08585_;
  assign _08588_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [7] : \MSYNC_1r1w.synth.nz.mem[356] [7];
  assign _08589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [7] : \MSYNC_1r1w.synth.nz.mem[358] [7];
  assign _08590_ = \bapg_rd.w_ptr_r [1] ? _08589_ : _08588_;
  assign _08591_ = \bapg_rd.w_ptr_r [2] ? _08590_ : _08587_;
  assign _08592_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [7] : \MSYNC_1r1w.synth.nz.mem[360] [7];
  assign _08593_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [7] : \MSYNC_1r1w.synth.nz.mem[362] [7];
  assign _08594_ = \bapg_rd.w_ptr_r [1] ? _08593_ : _08592_;
  assign _08595_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [7] : \MSYNC_1r1w.synth.nz.mem[364] [7];
  assign _08596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [7] : \MSYNC_1r1w.synth.nz.mem[366] [7];
  assign _08597_ = \bapg_rd.w_ptr_r [1] ? _08596_ : _08595_;
  assign _08598_ = \bapg_rd.w_ptr_r [2] ? _08597_ : _08594_;
  assign _08599_ = \bapg_rd.w_ptr_r [3] ? _08598_ : _08591_;
  assign _08600_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [7] : \MSYNC_1r1w.synth.nz.mem[368] [7];
  assign _08601_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [7] : \MSYNC_1r1w.synth.nz.mem[370] [7];
  assign _08602_ = \bapg_rd.w_ptr_r [1] ? _08601_ : _08600_;
  assign _08603_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [7] : \MSYNC_1r1w.synth.nz.mem[372] [7];
  assign _08604_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [7] : \MSYNC_1r1w.synth.nz.mem[374] [7];
  assign _08605_ = \bapg_rd.w_ptr_r [1] ? _08604_ : _08603_;
  assign _08606_ = \bapg_rd.w_ptr_r [2] ? _08605_ : _08602_;
  assign _08607_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [7] : \MSYNC_1r1w.synth.nz.mem[376] [7];
  assign _08608_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [7] : \MSYNC_1r1w.synth.nz.mem[378] [7];
  assign _08609_ = \bapg_rd.w_ptr_r [1] ? _08608_ : _08607_;
  assign _08610_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [7] : \MSYNC_1r1w.synth.nz.mem[380] [7];
  assign _08611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [7] : \MSYNC_1r1w.synth.nz.mem[382] [7];
  assign _08612_ = \bapg_rd.w_ptr_r [1] ? _08611_ : _08610_;
  assign _08613_ = \bapg_rd.w_ptr_r [2] ? _08612_ : _08609_;
  assign _08614_ = \bapg_rd.w_ptr_r [3] ? _08613_ : _08606_;
  assign _08615_ = \bapg_rd.w_ptr_r [4] ? _08614_ : _08599_;
  assign _08616_ = \bapg_rd.w_ptr_r [5] ? _08615_ : _08584_;
  assign _08617_ = \bapg_rd.w_ptr_r [6] ? _08616_ : _08553_;
  assign _08618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [7] : \MSYNC_1r1w.synth.nz.mem[384] [7];
  assign _08619_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [7] : \MSYNC_1r1w.synth.nz.mem[386] [7];
  assign _08620_ = \bapg_rd.w_ptr_r [1] ? _08619_ : _08618_;
  assign _08621_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [7] : \MSYNC_1r1w.synth.nz.mem[388] [7];
  assign _08622_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [7] : \MSYNC_1r1w.synth.nz.mem[390] [7];
  assign _08623_ = \bapg_rd.w_ptr_r [1] ? _08622_ : _08621_;
  assign _08624_ = \bapg_rd.w_ptr_r [2] ? _08623_ : _08620_;
  assign _08625_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [7] : \MSYNC_1r1w.synth.nz.mem[392] [7];
  assign _08626_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [7] : \MSYNC_1r1w.synth.nz.mem[394] [7];
  assign _08627_ = \bapg_rd.w_ptr_r [1] ? _08626_ : _08625_;
  assign _08628_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [7] : \MSYNC_1r1w.synth.nz.mem[396] [7];
  assign _08629_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [7] : \MSYNC_1r1w.synth.nz.mem[398] [7];
  assign _08630_ = \bapg_rd.w_ptr_r [1] ? _08629_ : _08628_;
  assign _08631_ = \bapg_rd.w_ptr_r [2] ? _08630_ : _08627_;
  assign _08632_ = \bapg_rd.w_ptr_r [3] ? _08631_ : _08624_;
  assign _08633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [7] : \MSYNC_1r1w.synth.nz.mem[400] [7];
  assign _08634_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [7] : \MSYNC_1r1w.synth.nz.mem[402] [7];
  assign _08635_ = \bapg_rd.w_ptr_r [1] ? _08634_ : _08633_;
  assign _08636_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [7] : \MSYNC_1r1w.synth.nz.mem[404] [7];
  assign _08637_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [7] : \MSYNC_1r1w.synth.nz.mem[406] [7];
  assign _08638_ = \bapg_rd.w_ptr_r [1] ? _08637_ : _08636_;
  assign _08639_ = \bapg_rd.w_ptr_r [2] ? _08638_ : _08635_;
  assign _08640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [7] : \MSYNC_1r1w.synth.nz.mem[408] [7];
  assign _08641_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [7] : \MSYNC_1r1w.synth.nz.mem[410] [7];
  assign _08642_ = \bapg_rd.w_ptr_r [1] ? _08641_ : _08640_;
  assign _08643_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [7] : \MSYNC_1r1w.synth.nz.mem[412] [7];
  assign _08644_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [7] : \MSYNC_1r1w.synth.nz.mem[414] [7];
  assign _08645_ = \bapg_rd.w_ptr_r [1] ? _08644_ : _08643_;
  assign _08646_ = \bapg_rd.w_ptr_r [2] ? _08645_ : _08642_;
  assign _08647_ = \bapg_rd.w_ptr_r [3] ? _08646_ : _08639_;
  assign _08648_ = \bapg_rd.w_ptr_r [4] ? _08647_ : _08632_;
  assign _08649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [7] : \MSYNC_1r1w.synth.nz.mem[416] [7];
  assign _08650_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [7] : \MSYNC_1r1w.synth.nz.mem[418] [7];
  assign _08651_ = \bapg_rd.w_ptr_r [1] ? _08650_ : _08649_;
  assign _08652_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [7] : \MSYNC_1r1w.synth.nz.mem[420] [7];
  assign _08653_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [7] : \MSYNC_1r1w.synth.nz.mem[422] [7];
  assign _08654_ = \bapg_rd.w_ptr_r [1] ? _08653_ : _08652_;
  assign _08655_ = \bapg_rd.w_ptr_r [2] ? _08654_ : _08651_;
  assign _08656_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [7] : \MSYNC_1r1w.synth.nz.mem[424] [7];
  assign _08657_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [7] : \MSYNC_1r1w.synth.nz.mem[426] [7];
  assign _08658_ = \bapg_rd.w_ptr_r [1] ? _08657_ : _08656_;
  assign _08659_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [7] : \MSYNC_1r1w.synth.nz.mem[428] [7];
  assign _08660_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [7] : \MSYNC_1r1w.synth.nz.mem[430] [7];
  assign _08661_ = \bapg_rd.w_ptr_r [1] ? _08660_ : _08659_;
  assign _08662_ = \bapg_rd.w_ptr_r [2] ? _08661_ : _08658_;
  assign _08663_ = \bapg_rd.w_ptr_r [3] ? _08662_ : _08655_;
  assign _08664_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [7] : \MSYNC_1r1w.synth.nz.mem[432] [7];
  assign _08665_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [7] : \MSYNC_1r1w.synth.nz.mem[434] [7];
  assign _08666_ = \bapg_rd.w_ptr_r [1] ? _08665_ : _08664_;
  assign _08667_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [7] : \MSYNC_1r1w.synth.nz.mem[436] [7];
  assign _08668_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [7] : \MSYNC_1r1w.synth.nz.mem[438] [7];
  assign _08669_ = \bapg_rd.w_ptr_r [1] ? _08668_ : _08667_;
  assign _08670_ = \bapg_rd.w_ptr_r [2] ? _08669_ : _08666_;
  assign _08671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [7] : \MSYNC_1r1w.synth.nz.mem[440] [7];
  assign _08672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [7] : \MSYNC_1r1w.synth.nz.mem[442] [7];
  assign _08673_ = \bapg_rd.w_ptr_r [1] ? _08672_ : _08671_;
  assign _08674_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [7] : \MSYNC_1r1w.synth.nz.mem[444] [7];
  assign _08675_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [7] : \MSYNC_1r1w.synth.nz.mem[446] [7];
  assign _08676_ = \bapg_rd.w_ptr_r [1] ? _08675_ : _08674_;
  assign _08677_ = \bapg_rd.w_ptr_r [2] ? _08676_ : _08673_;
  assign _08678_ = \bapg_rd.w_ptr_r [3] ? _08677_ : _08670_;
  assign _08679_ = \bapg_rd.w_ptr_r [4] ? _08678_ : _08663_;
  assign _08680_ = \bapg_rd.w_ptr_r [5] ? _08679_ : _08648_;
  assign _08681_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [7] : \MSYNC_1r1w.synth.nz.mem[448] [7];
  assign _08682_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [7] : \MSYNC_1r1w.synth.nz.mem[450] [7];
  assign _08683_ = \bapg_rd.w_ptr_r [1] ? _08682_ : _08681_;
  assign _08684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [7] : \MSYNC_1r1w.synth.nz.mem[452] [7];
  assign _08685_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [7] : \MSYNC_1r1w.synth.nz.mem[454] [7];
  assign _08686_ = \bapg_rd.w_ptr_r [1] ? _08685_ : _08684_;
  assign _08687_ = \bapg_rd.w_ptr_r [2] ? _08686_ : _08683_;
  assign _08688_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [7] : \MSYNC_1r1w.synth.nz.mem[456] [7];
  assign _08689_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [7] : \MSYNC_1r1w.synth.nz.mem[458] [7];
  assign _08690_ = \bapg_rd.w_ptr_r [1] ? _08689_ : _08688_;
  assign _08691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [7] : \MSYNC_1r1w.synth.nz.mem[460] [7];
  assign _08692_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [7] : \MSYNC_1r1w.synth.nz.mem[462] [7];
  assign _08693_ = \bapg_rd.w_ptr_r [1] ? _08692_ : _08691_;
  assign _08694_ = \bapg_rd.w_ptr_r [2] ? _08693_ : _08690_;
  assign _08695_ = \bapg_rd.w_ptr_r [3] ? _08694_ : _08687_;
  assign _08696_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [7] : \MSYNC_1r1w.synth.nz.mem[464] [7];
  assign _08697_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [7] : \MSYNC_1r1w.synth.nz.mem[466] [7];
  assign _08698_ = \bapg_rd.w_ptr_r [1] ? _08697_ : _08696_;
  assign _08699_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [7] : \MSYNC_1r1w.synth.nz.mem[468] [7];
  assign _08700_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [7] : \MSYNC_1r1w.synth.nz.mem[470] [7];
  assign _08701_ = \bapg_rd.w_ptr_r [1] ? _08700_ : _08699_;
  assign _08702_ = \bapg_rd.w_ptr_r [2] ? _08701_ : _08698_;
  assign _08703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [7] : \MSYNC_1r1w.synth.nz.mem[472] [7];
  assign _08704_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [7] : \MSYNC_1r1w.synth.nz.mem[474] [7];
  assign _08705_ = \bapg_rd.w_ptr_r [1] ? _08704_ : _08703_;
  assign _08706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [7] : \MSYNC_1r1w.synth.nz.mem[476] [7];
  assign _08707_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [7] : \MSYNC_1r1w.synth.nz.mem[478] [7];
  assign _08708_ = \bapg_rd.w_ptr_r [1] ? _08707_ : _08706_;
  assign _08709_ = \bapg_rd.w_ptr_r [2] ? _08708_ : _08705_;
  assign _08710_ = \bapg_rd.w_ptr_r [3] ? _08709_ : _08702_;
  assign _08711_ = \bapg_rd.w_ptr_r [4] ? _08710_ : _08695_;
  assign _08712_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [7] : \MSYNC_1r1w.synth.nz.mem[480] [7];
  assign _08713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [7] : \MSYNC_1r1w.synth.nz.mem[482] [7];
  assign _08714_ = \bapg_rd.w_ptr_r [1] ? _08713_ : _08712_;
  assign _08715_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [7] : \MSYNC_1r1w.synth.nz.mem[484] [7];
  assign _08716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [7] : \MSYNC_1r1w.synth.nz.mem[486] [7];
  assign _08717_ = \bapg_rd.w_ptr_r [1] ? _08716_ : _08715_;
  assign _08718_ = \bapg_rd.w_ptr_r [2] ? _08717_ : _08714_;
  assign _08719_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [7] : \MSYNC_1r1w.synth.nz.mem[488] [7];
  assign _08720_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [7] : \MSYNC_1r1w.synth.nz.mem[490] [7];
  assign _08721_ = \bapg_rd.w_ptr_r [1] ? _08720_ : _08719_;
  assign _08722_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [7] : \MSYNC_1r1w.synth.nz.mem[492] [7];
  assign _08723_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [7] : \MSYNC_1r1w.synth.nz.mem[494] [7];
  assign _08724_ = \bapg_rd.w_ptr_r [1] ? _08723_ : _08722_;
  assign _08725_ = \bapg_rd.w_ptr_r [2] ? _08724_ : _08721_;
  assign _08726_ = \bapg_rd.w_ptr_r [3] ? _08725_ : _08718_;
  assign _08727_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [7] : \MSYNC_1r1w.synth.nz.mem[496] [7];
  assign _08728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [7] : \MSYNC_1r1w.synth.nz.mem[498] [7];
  assign _08729_ = \bapg_rd.w_ptr_r [1] ? _08728_ : _08727_;
  assign _08730_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [7] : \MSYNC_1r1w.synth.nz.mem[500] [7];
  assign _08731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [7] : \MSYNC_1r1w.synth.nz.mem[502] [7];
  assign _08732_ = \bapg_rd.w_ptr_r [1] ? _08731_ : _08730_;
  assign _08733_ = \bapg_rd.w_ptr_r [2] ? _08732_ : _08729_;
  assign _08734_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [7] : \MSYNC_1r1w.synth.nz.mem[504] [7];
  assign _08735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [7] : \MSYNC_1r1w.synth.nz.mem[506] [7];
  assign _08736_ = \bapg_rd.w_ptr_r [1] ? _08735_ : _08734_;
  assign _08737_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [7] : \MSYNC_1r1w.synth.nz.mem[508] [7];
  assign _08738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [7] : \MSYNC_1r1w.synth.nz.mem[510] [7];
  assign _08739_ = \bapg_rd.w_ptr_r [1] ? _08738_ : _08737_;
  assign _08740_ = \bapg_rd.w_ptr_r [2] ? _08739_ : _08736_;
  assign _08741_ = \bapg_rd.w_ptr_r [3] ? _08740_ : _08733_;
  assign _08742_ = \bapg_rd.w_ptr_r [4] ? _08741_ : _08726_;
  assign _08743_ = \bapg_rd.w_ptr_r [5] ? _08742_ : _08711_;
  assign _08744_ = \bapg_rd.w_ptr_r [6] ? _08743_ : _08680_;
  assign _08745_ = \bapg_rd.w_ptr_r [7] ? _08744_ : _08617_;
  assign _08746_ = \bapg_rd.w_ptr_r [8] ? _08745_ : _08490_;
  assign _08747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [7] : \MSYNC_1r1w.synth.nz.mem[512] [7];
  assign _08748_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [7] : \MSYNC_1r1w.synth.nz.mem[514] [7];
  assign _08749_ = \bapg_rd.w_ptr_r [1] ? _08748_ : _08747_;
  assign _08750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [7] : \MSYNC_1r1w.synth.nz.mem[516] [7];
  assign _08751_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [7] : \MSYNC_1r1w.synth.nz.mem[518] [7];
  assign _08752_ = \bapg_rd.w_ptr_r [1] ? _08751_ : _08750_;
  assign _08753_ = \bapg_rd.w_ptr_r [2] ? _08752_ : _08749_;
  assign _08754_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [7] : \MSYNC_1r1w.synth.nz.mem[520] [7];
  assign _08755_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [7] : \MSYNC_1r1w.synth.nz.mem[522] [7];
  assign _08756_ = \bapg_rd.w_ptr_r [1] ? _08755_ : _08754_;
  assign _08757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [7] : \MSYNC_1r1w.synth.nz.mem[524] [7];
  assign _08758_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [7] : \MSYNC_1r1w.synth.nz.mem[526] [7];
  assign _08759_ = \bapg_rd.w_ptr_r [1] ? _08758_ : _08757_;
  assign _08760_ = \bapg_rd.w_ptr_r [2] ? _08759_ : _08756_;
  assign _08761_ = \bapg_rd.w_ptr_r [3] ? _08760_ : _08753_;
  assign _08762_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [7] : \MSYNC_1r1w.synth.nz.mem[528] [7];
  assign _08763_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [7] : \MSYNC_1r1w.synth.nz.mem[530] [7];
  assign _08764_ = \bapg_rd.w_ptr_r [1] ? _08763_ : _08762_;
  assign _08765_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [7] : \MSYNC_1r1w.synth.nz.mem[532] [7];
  assign _08766_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [7] : \MSYNC_1r1w.synth.nz.mem[534] [7];
  assign _08767_ = \bapg_rd.w_ptr_r [1] ? _08766_ : _08765_;
  assign _08768_ = \bapg_rd.w_ptr_r [2] ? _08767_ : _08764_;
  assign _08769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [7] : \MSYNC_1r1w.synth.nz.mem[536] [7];
  assign _08770_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [7] : \MSYNC_1r1w.synth.nz.mem[538] [7];
  assign _08771_ = \bapg_rd.w_ptr_r [1] ? _08770_ : _08769_;
  assign _08772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [7] : \MSYNC_1r1w.synth.nz.mem[540] [7];
  assign _08773_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [7] : \MSYNC_1r1w.synth.nz.mem[542] [7];
  assign _08774_ = \bapg_rd.w_ptr_r [1] ? _08773_ : _08772_;
  assign _08775_ = \bapg_rd.w_ptr_r [2] ? _08774_ : _08771_;
  assign _08776_ = \bapg_rd.w_ptr_r [3] ? _08775_ : _08768_;
  assign _08777_ = \bapg_rd.w_ptr_r [4] ? _08776_ : _08761_;
  assign _08778_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [7] : \MSYNC_1r1w.synth.nz.mem[544] [7];
  assign _08779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [7] : \MSYNC_1r1w.synth.nz.mem[546] [7];
  assign _08780_ = \bapg_rd.w_ptr_r [1] ? _08779_ : _08778_;
  assign _08781_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [7] : \MSYNC_1r1w.synth.nz.mem[548] [7];
  assign _08782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [7] : \MSYNC_1r1w.synth.nz.mem[550] [7];
  assign _08783_ = \bapg_rd.w_ptr_r [1] ? _08782_ : _08781_;
  assign _08784_ = \bapg_rd.w_ptr_r [2] ? _08783_ : _08780_;
  assign _08785_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [7] : \MSYNC_1r1w.synth.nz.mem[552] [7];
  assign _08786_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [7] : \MSYNC_1r1w.synth.nz.mem[554] [7];
  assign _08787_ = \bapg_rd.w_ptr_r [1] ? _08786_ : _08785_;
  assign _08788_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [7] : \MSYNC_1r1w.synth.nz.mem[556] [7];
  assign _08789_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [7] : \MSYNC_1r1w.synth.nz.mem[558] [7];
  assign _08790_ = \bapg_rd.w_ptr_r [1] ? _08789_ : _08788_;
  assign _08791_ = \bapg_rd.w_ptr_r [2] ? _08790_ : _08787_;
  assign _08792_ = \bapg_rd.w_ptr_r [3] ? _08791_ : _08784_;
  assign _08793_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [7] : \MSYNC_1r1w.synth.nz.mem[560] [7];
  assign _08794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [7] : \MSYNC_1r1w.synth.nz.mem[562] [7];
  assign _08795_ = \bapg_rd.w_ptr_r [1] ? _08794_ : _08793_;
  assign _08796_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [7] : \MSYNC_1r1w.synth.nz.mem[564] [7];
  assign _08797_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [7] : \MSYNC_1r1w.synth.nz.mem[566] [7];
  assign _08798_ = \bapg_rd.w_ptr_r [1] ? _08797_ : _08796_;
  assign _08799_ = \bapg_rd.w_ptr_r [2] ? _08798_ : _08795_;
  assign _08800_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [7] : \MSYNC_1r1w.synth.nz.mem[568] [7];
  assign _08801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [7] : \MSYNC_1r1w.synth.nz.mem[570] [7];
  assign _08802_ = \bapg_rd.w_ptr_r [1] ? _08801_ : _08800_;
  assign _08803_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [7] : \MSYNC_1r1w.synth.nz.mem[572] [7];
  assign _08804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [7] : \MSYNC_1r1w.synth.nz.mem[574] [7];
  assign _08805_ = \bapg_rd.w_ptr_r [1] ? _08804_ : _08803_;
  assign _08806_ = \bapg_rd.w_ptr_r [2] ? _08805_ : _08802_;
  assign _08807_ = \bapg_rd.w_ptr_r [3] ? _08806_ : _08799_;
  assign _08808_ = \bapg_rd.w_ptr_r [4] ? _08807_ : _08792_;
  assign _08809_ = \bapg_rd.w_ptr_r [5] ? _08808_ : _08777_;
  assign _08810_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [7] : \MSYNC_1r1w.synth.nz.mem[576] [7];
  assign _08811_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [7] : \MSYNC_1r1w.synth.nz.mem[578] [7];
  assign _08812_ = \bapg_rd.w_ptr_r [1] ? _08811_ : _08810_;
  assign _08813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [7] : \MSYNC_1r1w.synth.nz.mem[580] [7];
  assign _08814_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [7] : \MSYNC_1r1w.synth.nz.mem[582] [7];
  assign _08815_ = \bapg_rd.w_ptr_r [1] ? _08814_ : _08813_;
  assign _08816_ = \bapg_rd.w_ptr_r [2] ? _08815_ : _08812_;
  assign _08817_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [7] : \MSYNC_1r1w.synth.nz.mem[584] [7];
  assign _08818_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [7] : \MSYNC_1r1w.synth.nz.mem[586] [7];
  assign _08819_ = \bapg_rd.w_ptr_r [1] ? _08818_ : _08817_;
  assign _08820_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [7] : \MSYNC_1r1w.synth.nz.mem[588] [7];
  assign _08821_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [7] : \MSYNC_1r1w.synth.nz.mem[590] [7];
  assign _08822_ = \bapg_rd.w_ptr_r [1] ? _08821_ : _08820_;
  assign _08823_ = \bapg_rd.w_ptr_r [2] ? _08822_ : _08819_;
  assign _08824_ = \bapg_rd.w_ptr_r [3] ? _08823_ : _08816_;
  assign _08825_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [7] : \MSYNC_1r1w.synth.nz.mem[592] [7];
  assign _08826_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [7] : \MSYNC_1r1w.synth.nz.mem[594] [7];
  assign _08827_ = \bapg_rd.w_ptr_r [1] ? _08826_ : _08825_;
  assign _08828_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [7] : \MSYNC_1r1w.synth.nz.mem[596] [7];
  assign _08829_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [7] : \MSYNC_1r1w.synth.nz.mem[598] [7];
  assign _08830_ = \bapg_rd.w_ptr_r [1] ? _08829_ : _08828_;
  assign _08831_ = \bapg_rd.w_ptr_r [2] ? _08830_ : _08827_;
  assign _08832_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [7] : \MSYNC_1r1w.synth.nz.mem[600] [7];
  assign _08833_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [7] : \MSYNC_1r1w.synth.nz.mem[602] [7];
  assign _08834_ = \bapg_rd.w_ptr_r [1] ? _08833_ : _08832_;
  assign _08835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [7] : \MSYNC_1r1w.synth.nz.mem[604] [7];
  assign _08836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [7] : \MSYNC_1r1w.synth.nz.mem[606] [7];
  assign _08837_ = \bapg_rd.w_ptr_r [1] ? _08836_ : _08835_;
  assign _08838_ = \bapg_rd.w_ptr_r [2] ? _08837_ : _08834_;
  assign _08839_ = \bapg_rd.w_ptr_r [3] ? _08838_ : _08831_;
  assign _08840_ = \bapg_rd.w_ptr_r [4] ? _08839_ : _08824_;
  assign _08841_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [7] : \MSYNC_1r1w.synth.nz.mem[608] [7];
  assign _08842_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [7] : \MSYNC_1r1w.synth.nz.mem[610] [7];
  assign _08843_ = \bapg_rd.w_ptr_r [1] ? _08842_ : _08841_;
  assign _08844_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [7] : \MSYNC_1r1w.synth.nz.mem[612] [7];
  assign _08845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [7] : \MSYNC_1r1w.synth.nz.mem[614] [7];
  assign _08846_ = \bapg_rd.w_ptr_r [1] ? _08845_ : _08844_;
  assign _08847_ = \bapg_rd.w_ptr_r [2] ? _08846_ : _08843_;
  assign _08848_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [7] : \MSYNC_1r1w.synth.nz.mem[616] [7];
  assign _08849_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [7] : \MSYNC_1r1w.synth.nz.mem[618] [7];
  assign _08850_ = \bapg_rd.w_ptr_r [1] ? _08849_ : _08848_;
  assign _08851_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [7] : \MSYNC_1r1w.synth.nz.mem[620] [7];
  assign _08852_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [7] : \MSYNC_1r1w.synth.nz.mem[622] [7];
  assign _08853_ = \bapg_rd.w_ptr_r [1] ? _08852_ : _08851_;
  assign _08854_ = \bapg_rd.w_ptr_r [2] ? _08853_ : _08850_;
  assign _08855_ = \bapg_rd.w_ptr_r [3] ? _08854_ : _08847_;
  assign _08856_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [7] : \MSYNC_1r1w.synth.nz.mem[624] [7];
  assign _08857_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [7] : \MSYNC_1r1w.synth.nz.mem[626] [7];
  assign _08858_ = \bapg_rd.w_ptr_r [1] ? _08857_ : _08856_;
  assign _08859_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [7] : \MSYNC_1r1w.synth.nz.mem[628] [7];
  assign _08860_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [7] : \MSYNC_1r1w.synth.nz.mem[630] [7];
  assign _08861_ = \bapg_rd.w_ptr_r [1] ? _08860_ : _08859_;
  assign _08862_ = \bapg_rd.w_ptr_r [2] ? _08861_ : _08858_;
  assign _08863_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [7] : \MSYNC_1r1w.synth.nz.mem[632] [7];
  assign _08864_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [7] : \MSYNC_1r1w.synth.nz.mem[634] [7];
  assign _08865_ = \bapg_rd.w_ptr_r [1] ? _08864_ : _08863_;
  assign _08866_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [7] : \MSYNC_1r1w.synth.nz.mem[636] [7];
  assign _08867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [7] : \MSYNC_1r1w.synth.nz.mem[638] [7];
  assign _08868_ = \bapg_rd.w_ptr_r [1] ? _08867_ : _08866_;
  assign _08869_ = \bapg_rd.w_ptr_r [2] ? _08868_ : _08865_;
  assign _08870_ = \bapg_rd.w_ptr_r [3] ? _08869_ : _08862_;
  assign _08871_ = \bapg_rd.w_ptr_r [4] ? _08870_ : _08855_;
  assign _08872_ = \bapg_rd.w_ptr_r [5] ? _08871_ : _08840_;
  assign _08873_ = \bapg_rd.w_ptr_r [6] ? _08872_ : _08809_;
  assign _08874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [7] : \MSYNC_1r1w.synth.nz.mem[640] [7];
  assign _08875_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [7] : \MSYNC_1r1w.synth.nz.mem[642] [7];
  assign _08876_ = \bapg_rd.w_ptr_r [1] ? _08875_ : _08874_;
  assign _08877_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [7] : \MSYNC_1r1w.synth.nz.mem[644] [7];
  assign _08878_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [7] : \MSYNC_1r1w.synth.nz.mem[646] [7];
  assign _08879_ = \bapg_rd.w_ptr_r [1] ? _08878_ : _08877_;
  assign _08880_ = \bapg_rd.w_ptr_r [2] ? _08879_ : _08876_;
  assign _08881_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [7] : \MSYNC_1r1w.synth.nz.mem[648] [7];
  assign _08882_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [7] : \MSYNC_1r1w.synth.nz.mem[650] [7];
  assign _08883_ = \bapg_rd.w_ptr_r [1] ? _08882_ : _08881_;
  assign _08884_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [7] : \MSYNC_1r1w.synth.nz.mem[652] [7];
  assign _08885_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [7] : \MSYNC_1r1w.synth.nz.mem[654] [7];
  assign _08886_ = \bapg_rd.w_ptr_r [1] ? _08885_ : _08884_;
  assign _08887_ = \bapg_rd.w_ptr_r [2] ? _08886_ : _08883_;
  assign _08888_ = \bapg_rd.w_ptr_r [3] ? _08887_ : _08880_;
  assign _08889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [7] : \MSYNC_1r1w.synth.nz.mem[656] [7];
  assign _08890_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [7] : \MSYNC_1r1w.synth.nz.mem[658] [7];
  assign _08891_ = \bapg_rd.w_ptr_r [1] ? _08890_ : _08889_;
  assign _08892_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [7] : \MSYNC_1r1w.synth.nz.mem[660] [7];
  assign _08893_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [7] : \MSYNC_1r1w.synth.nz.mem[662] [7];
  assign _08894_ = \bapg_rd.w_ptr_r [1] ? _08893_ : _08892_;
  assign _08895_ = \bapg_rd.w_ptr_r [2] ? _08894_ : _08891_;
  assign _08896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [7] : \MSYNC_1r1w.synth.nz.mem[664] [7];
  assign _08897_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [7] : \MSYNC_1r1w.synth.nz.mem[666] [7];
  assign _08898_ = \bapg_rd.w_ptr_r [1] ? _08897_ : _08896_;
  assign _08899_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [7] : \MSYNC_1r1w.synth.nz.mem[668] [7];
  assign _08900_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [7] : \MSYNC_1r1w.synth.nz.mem[670] [7];
  assign _08901_ = \bapg_rd.w_ptr_r [1] ? _08900_ : _08899_;
  assign _08902_ = \bapg_rd.w_ptr_r [2] ? _08901_ : _08898_;
  assign _08903_ = \bapg_rd.w_ptr_r [3] ? _08902_ : _08895_;
  assign _08904_ = \bapg_rd.w_ptr_r [4] ? _08903_ : _08888_;
  assign _08905_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [7] : \MSYNC_1r1w.synth.nz.mem[672] [7];
  assign _08906_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [7] : \MSYNC_1r1w.synth.nz.mem[674] [7];
  assign _08907_ = \bapg_rd.w_ptr_r [1] ? _08906_ : _08905_;
  assign _08908_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [7] : \MSYNC_1r1w.synth.nz.mem[676] [7];
  assign _08909_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [7] : \MSYNC_1r1w.synth.nz.mem[678] [7];
  assign _08910_ = \bapg_rd.w_ptr_r [1] ? _08909_ : _08908_;
  assign _08911_ = \bapg_rd.w_ptr_r [2] ? _08910_ : _08907_;
  assign _08912_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [7] : \MSYNC_1r1w.synth.nz.mem[680] [7];
  assign _08913_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [7] : \MSYNC_1r1w.synth.nz.mem[682] [7];
  assign _08914_ = \bapg_rd.w_ptr_r [1] ? _08913_ : _08912_;
  assign _08915_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [7] : \MSYNC_1r1w.synth.nz.mem[684] [7];
  assign _08916_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [7] : \MSYNC_1r1w.synth.nz.mem[686] [7];
  assign _08917_ = \bapg_rd.w_ptr_r [1] ? _08916_ : _08915_;
  assign _08918_ = \bapg_rd.w_ptr_r [2] ? _08917_ : _08914_;
  assign _08919_ = \bapg_rd.w_ptr_r [3] ? _08918_ : _08911_;
  assign _08920_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [7] : \MSYNC_1r1w.synth.nz.mem[688] [7];
  assign _08921_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [7] : \MSYNC_1r1w.synth.nz.mem[690] [7];
  assign _08922_ = \bapg_rd.w_ptr_r [1] ? _08921_ : _08920_;
  assign _08923_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [7] : \MSYNC_1r1w.synth.nz.mem[692] [7];
  assign _08924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [7] : \MSYNC_1r1w.synth.nz.mem[694] [7];
  assign _08925_ = \bapg_rd.w_ptr_r [1] ? _08924_ : _08923_;
  assign _08926_ = \bapg_rd.w_ptr_r [2] ? _08925_ : _08922_;
  assign _08927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [7] : \MSYNC_1r1w.synth.nz.mem[696] [7];
  assign _08928_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [7] : \MSYNC_1r1w.synth.nz.mem[698] [7];
  assign _08929_ = \bapg_rd.w_ptr_r [1] ? _08928_ : _08927_;
  assign _08930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [7] : \MSYNC_1r1w.synth.nz.mem[700] [7];
  assign _08931_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [7] : \MSYNC_1r1w.synth.nz.mem[702] [7];
  assign _08932_ = \bapg_rd.w_ptr_r [1] ? _08931_ : _08930_;
  assign _08933_ = \bapg_rd.w_ptr_r [2] ? _08932_ : _08929_;
  assign _08934_ = \bapg_rd.w_ptr_r [3] ? _08933_ : _08926_;
  assign _08935_ = \bapg_rd.w_ptr_r [4] ? _08934_ : _08919_;
  assign _08936_ = \bapg_rd.w_ptr_r [5] ? _08935_ : _08904_;
  assign _08937_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [7] : \MSYNC_1r1w.synth.nz.mem[704] [7];
  assign _08938_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [7] : \MSYNC_1r1w.synth.nz.mem[706] [7];
  assign _08939_ = \bapg_rd.w_ptr_r [1] ? _08938_ : _08937_;
  assign _08940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [7] : \MSYNC_1r1w.synth.nz.mem[708] [7];
  assign _08941_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [7] : \MSYNC_1r1w.synth.nz.mem[710] [7];
  assign _08942_ = \bapg_rd.w_ptr_r [1] ? _08941_ : _08940_;
  assign _08943_ = \bapg_rd.w_ptr_r [2] ? _08942_ : _08939_;
  assign _08944_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [7] : \MSYNC_1r1w.synth.nz.mem[712] [7];
  assign _08945_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [7] : \MSYNC_1r1w.synth.nz.mem[714] [7];
  assign _08946_ = \bapg_rd.w_ptr_r [1] ? _08945_ : _08944_;
  assign _08947_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [7] : \MSYNC_1r1w.synth.nz.mem[716] [7];
  assign _08948_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [7] : \MSYNC_1r1w.synth.nz.mem[718] [7];
  assign _08949_ = \bapg_rd.w_ptr_r [1] ? _08948_ : _08947_;
  assign _08950_ = \bapg_rd.w_ptr_r [2] ? _08949_ : _08946_;
  assign _08951_ = \bapg_rd.w_ptr_r [3] ? _08950_ : _08943_;
  assign _08952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [7] : \MSYNC_1r1w.synth.nz.mem[720] [7];
  assign _08953_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [7] : \MSYNC_1r1w.synth.nz.mem[722] [7];
  assign _08954_ = \bapg_rd.w_ptr_r [1] ? _08953_ : _08952_;
  assign _08955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [7] : \MSYNC_1r1w.synth.nz.mem[724] [7];
  assign _08956_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [7] : \MSYNC_1r1w.synth.nz.mem[726] [7];
  assign _08957_ = \bapg_rd.w_ptr_r [1] ? _08956_ : _08955_;
  assign _08958_ = \bapg_rd.w_ptr_r [2] ? _08957_ : _08954_;
  assign _08959_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [7] : \MSYNC_1r1w.synth.nz.mem[728] [7];
  assign _08960_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [7] : \MSYNC_1r1w.synth.nz.mem[730] [7];
  assign _08961_ = \bapg_rd.w_ptr_r [1] ? _08960_ : _08959_;
  assign _08962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [7] : \MSYNC_1r1w.synth.nz.mem[732] [7];
  assign _08963_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [7] : \MSYNC_1r1w.synth.nz.mem[734] [7];
  assign _08964_ = \bapg_rd.w_ptr_r [1] ? _08963_ : _08962_;
  assign _08965_ = \bapg_rd.w_ptr_r [2] ? _08964_ : _08961_;
  assign _08966_ = \bapg_rd.w_ptr_r [3] ? _08965_ : _08958_;
  assign _08967_ = \bapg_rd.w_ptr_r [4] ? _08966_ : _08951_;
  assign _08968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [7] : \MSYNC_1r1w.synth.nz.mem[736] [7];
  assign _08969_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [7] : \MSYNC_1r1w.synth.nz.mem[738] [7];
  assign _08970_ = \bapg_rd.w_ptr_r [1] ? _08969_ : _08968_;
  assign _08971_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [7] : \MSYNC_1r1w.synth.nz.mem[740] [7];
  assign _08972_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [7] : \MSYNC_1r1w.synth.nz.mem[742] [7];
  assign _08973_ = \bapg_rd.w_ptr_r [1] ? _08972_ : _08971_;
  assign _08974_ = \bapg_rd.w_ptr_r [2] ? _08973_ : _08970_;
  assign _08975_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [7] : \MSYNC_1r1w.synth.nz.mem[744] [7];
  assign _08976_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [7] : \MSYNC_1r1w.synth.nz.mem[746] [7];
  assign _08977_ = \bapg_rd.w_ptr_r [1] ? _08976_ : _08975_;
  assign _08978_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [7] : \MSYNC_1r1w.synth.nz.mem[748] [7];
  assign _08979_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [7] : \MSYNC_1r1w.synth.nz.mem[750] [7];
  assign _08980_ = \bapg_rd.w_ptr_r [1] ? _08979_ : _08978_;
  assign _08981_ = \bapg_rd.w_ptr_r [2] ? _08980_ : _08977_;
  assign _08982_ = \bapg_rd.w_ptr_r [3] ? _08981_ : _08974_;
  assign _08983_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [7] : \MSYNC_1r1w.synth.nz.mem[752] [7];
  assign _08984_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [7] : \MSYNC_1r1w.synth.nz.mem[754] [7];
  assign _08985_ = \bapg_rd.w_ptr_r [1] ? _08984_ : _08983_;
  assign _08986_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [7] : \MSYNC_1r1w.synth.nz.mem[756] [7];
  assign _08987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [7] : \MSYNC_1r1w.synth.nz.mem[758] [7];
  assign _08988_ = \bapg_rd.w_ptr_r [1] ? _08987_ : _08986_;
  assign _08989_ = \bapg_rd.w_ptr_r [2] ? _08988_ : _08985_;
  assign _08990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [7] : \MSYNC_1r1w.synth.nz.mem[760] [7];
  assign _08991_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [7] : \MSYNC_1r1w.synth.nz.mem[762] [7];
  assign _08992_ = \bapg_rd.w_ptr_r [1] ? _08991_ : _08990_;
  assign _08993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [7] : \MSYNC_1r1w.synth.nz.mem[764] [7];
  assign _08994_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [7] : \MSYNC_1r1w.synth.nz.mem[766] [7];
  assign _08995_ = \bapg_rd.w_ptr_r [1] ? _08994_ : _08993_;
  assign _08996_ = \bapg_rd.w_ptr_r [2] ? _08995_ : _08992_;
  assign _08997_ = \bapg_rd.w_ptr_r [3] ? _08996_ : _08989_;
  assign _08998_ = \bapg_rd.w_ptr_r [4] ? _08997_ : _08982_;
  assign _08999_ = \bapg_rd.w_ptr_r [5] ? _08998_ : _08967_;
  assign _09000_ = \bapg_rd.w_ptr_r [6] ? _08999_ : _08936_;
  assign _09001_ = \bapg_rd.w_ptr_r [7] ? _09000_ : _08873_;
  assign _09002_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [7] : \MSYNC_1r1w.synth.nz.mem[768] [7];
  assign _09003_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [7] : \MSYNC_1r1w.synth.nz.mem[770] [7];
  assign _09004_ = \bapg_rd.w_ptr_r [1] ? _09003_ : _09002_;
  assign _09005_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [7] : \MSYNC_1r1w.synth.nz.mem[772] [7];
  assign _09006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [7] : \MSYNC_1r1w.synth.nz.mem[774] [7];
  assign _09007_ = \bapg_rd.w_ptr_r [1] ? _09006_ : _09005_;
  assign _09008_ = \bapg_rd.w_ptr_r [2] ? _09007_ : _09004_;
  assign _09009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [7] : \MSYNC_1r1w.synth.nz.mem[776] [7];
  assign _09010_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [7] : \MSYNC_1r1w.synth.nz.mem[778] [7];
  assign _09011_ = \bapg_rd.w_ptr_r [1] ? _09010_ : _09009_;
  assign _09012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [7] : \MSYNC_1r1w.synth.nz.mem[780] [7];
  assign _09013_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [7] : \MSYNC_1r1w.synth.nz.mem[782] [7];
  assign _09014_ = \bapg_rd.w_ptr_r [1] ? _09013_ : _09012_;
  assign _09015_ = \bapg_rd.w_ptr_r [2] ? _09014_ : _09011_;
  assign _09016_ = \bapg_rd.w_ptr_r [3] ? _09015_ : _09008_;
  assign _09017_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [7] : \MSYNC_1r1w.synth.nz.mem[784] [7];
  assign _09018_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [7] : \MSYNC_1r1w.synth.nz.mem[786] [7];
  assign _09019_ = \bapg_rd.w_ptr_r [1] ? _09018_ : _09017_;
  assign _09020_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [7] : \MSYNC_1r1w.synth.nz.mem[788] [7];
  assign _09021_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [7] : \MSYNC_1r1w.synth.nz.mem[790] [7];
  assign _09022_ = \bapg_rd.w_ptr_r [1] ? _09021_ : _09020_;
  assign _09023_ = \bapg_rd.w_ptr_r [2] ? _09022_ : _09019_;
  assign _09024_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [7] : \MSYNC_1r1w.synth.nz.mem[792] [7];
  assign _09025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [7] : \MSYNC_1r1w.synth.nz.mem[794] [7];
  assign _09026_ = \bapg_rd.w_ptr_r [1] ? _09025_ : _09024_;
  assign _09027_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [7] : \MSYNC_1r1w.synth.nz.mem[796] [7];
  assign _09028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [7] : \MSYNC_1r1w.synth.nz.mem[798] [7];
  assign _09029_ = \bapg_rd.w_ptr_r [1] ? _09028_ : _09027_;
  assign _09030_ = \bapg_rd.w_ptr_r [2] ? _09029_ : _09026_;
  assign _09031_ = \bapg_rd.w_ptr_r [3] ? _09030_ : _09023_;
  assign _09032_ = \bapg_rd.w_ptr_r [4] ? _09031_ : _09016_;
  assign _09033_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [7] : \MSYNC_1r1w.synth.nz.mem[800] [7];
  assign _09034_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [7] : \MSYNC_1r1w.synth.nz.mem[802] [7];
  assign _09035_ = \bapg_rd.w_ptr_r [1] ? _09034_ : _09033_;
  assign _09036_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [7] : \MSYNC_1r1w.synth.nz.mem[804] [7];
  assign _09037_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [7] : \MSYNC_1r1w.synth.nz.mem[806] [7];
  assign _09038_ = \bapg_rd.w_ptr_r [1] ? _09037_ : _09036_;
  assign _09039_ = \bapg_rd.w_ptr_r [2] ? _09038_ : _09035_;
  assign _09040_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [7] : \MSYNC_1r1w.synth.nz.mem[808] [7];
  assign _09041_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [7] : \MSYNC_1r1w.synth.nz.mem[810] [7];
  assign _09042_ = \bapg_rd.w_ptr_r [1] ? _09041_ : _09040_;
  assign _09043_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [7] : \MSYNC_1r1w.synth.nz.mem[812] [7];
  assign _09044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [7] : \MSYNC_1r1w.synth.nz.mem[814] [7];
  assign _09045_ = \bapg_rd.w_ptr_r [1] ? _09044_ : _09043_;
  assign _09046_ = \bapg_rd.w_ptr_r [2] ? _09045_ : _09042_;
  assign _09047_ = \bapg_rd.w_ptr_r [3] ? _09046_ : _09039_;
  assign _09048_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [7] : \MSYNC_1r1w.synth.nz.mem[816] [7];
  assign _09049_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [7] : \MSYNC_1r1w.synth.nz.mem[818] [7];
  assign _09050_ = \bapg_rd.w_ptr_r [1] ? _09049_ : _09048_;
  assign _09051_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [7] : \MSYNC_1r1w.synth.nz.mem[820] [7];
  assign _09052_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [7] : \MSYNC_1r1w.synth.nz.mem[822] [7];
  assign _09053_ = \bapg_rd.w_ptr_r [1] ? _09052_ : _09051_;
  assign _09054_ = \bapg_rd.w_ptr_r [2] ? _09053_ : _09050_;
  assign _09055_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [7] : \MSYNC_1r1w.synth.nz.mem[824] [7];
  assign _09056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [7] : \MSYNC_1r1w.synth.nz.mem[826] [7];
  assign _09057_ = \bapg_rd.w_ptr_r [1] ? _09056_ : _09055_;
  assign _09058_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [7] : \MSYNC_1r1w.synth.nz.mem[828] [7];
  assign _09059_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [7] : \MSYNC_1r1w.synth.nz.mem[830] [7];
  assign _09060_ = \bapg_rd.w_ptr_r [1] ? _09059_ : _09058_;
  assign _09061_ = \bapg_rd.w_ptr_r [2] ? _09060_ : _09057_;
  assign _09062_ = \bapg_rd.w_ptr_r [3] ? _09061_ : _09054_;
  assign _09063_ = \bapg_rd.w_ptr_r [4] ? _09062_ : _09047_;
  assign _09064_ = \bapg_rd.w_ptr_r [5] ? _09063_ : _09032_;
  assign _09065_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [7] : \MSYNC_1r1w.synth.nz.mem[832] [7];
  assign _09066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [7] : \MSYNC_1r1w.synth.nz.mem[834] [7];
  assign _09067_ = \bapg_rd.w_ptr_r [1] ? _09066_ : _09065_;
  assign _09068_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [7] : \MSYNC_1r1w.synth.nz.mem[836] [7];
  assign _09069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [7] : \MSYNC_1r1w.synth.nz.mem[838] [7];
  assign _09070_ = \bapg_rd.w_ptr_r [1] ? _09069_ : _09068_;
  assign _09071_ = \bapg_rd.w_ptr_r [2] ? _09070_ : _09067_;
  assign _09072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [7] : \MSYNC_1r1w.synth.nz.mem[840] [7];
  assign _09073_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [7] : \MSYNC_1r1w.synth.nz.mem[842] [7];
  assign _09074_ = \bapg_rd.w_ptr_r [1] ? _09073_ : _09072_;
  assign _09075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [7] : \MSYNC_1r1w.synth.nz.mem[844] [7];
  assign _09076_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [7] : \MSYNC_1r1w.synth.nz.mem[846] [7];
  assign _09077_ = \bapg_rd.w_ptr_r [1] ? _09076_ : _09075_;
  assign _09078_ = \bapg_rd.w_ptr_r [2] ? _09077_ : _09074_;
  assign _09079_ = \bapg_rd.w_ptr_r [3] ? _09078_ : _09071_;
  assign _09080_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [7] : \MSYNC_1r1w.synth.nz.mem[848] [7];
  assign _09081_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [7] : \MSYNC_1r1w.synth.nz.mem[850] [7];
  assign _09082_ = \bapg_rd.w_ptr_r [1] ? _09081_ : _09080_;
  assign _09083_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [7] : \MSYNC_1r1w.synth.nz.mem[852] [7];
  assign _09084_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [7] : \MSYNC_1r1w.synth.nz.mem[854] [7];
  assign _09085_ = \bapg_rd.w_ptr_r [1] ? _09084_ : _09083_;
  assign _09086_ = \bapg_rd.w_ptr_r [2] ? _09085_ : _09082_;
  assign _09087_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [7] : \MSYNC_1r1w.synth.nz.mem[856] [7];
  assign _09088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [7] : \MSYNC_1r1w.synth.nz.mem[858] [7];
  assign _09089_ = \bapg_rd.w_ptr_r [1] ? _09088_ : _09087_;
  assign _09090_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [7] : \MSYNC_1r1w.synth.nz.mem[860] [7];
  assign _09091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [7] : \MSYNC_1r1w.synth.nz.mem[862] [7];
  assign _09092_ = \bapg_rd.w_ptr_r [1] ? _09091_ : _09090_;
  assign _09093_ = \bapg_rd.w_ptr_r [2] ? _09092_ : _09089_;
  assign _09094_ = \bapg_rd.w_ptr_r [3] ? _09093_ : _09086_;
  assign _09095_ = \bapg_rd.w_ptr_r [4] ? _09094_ : _09079_;
  assign _09096_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [7] : \MSYNC_1r1w.synth.nz.mem[864] [7];
  assign _09097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [7] : \MSYNC_1r1w.synth.nz.mem[866] [7];
  assign _09098_ = \bapg_rd.w_ptr_r [1] ? _09097_ : _09096_;
  assign _09099_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [7] : \MSYNC_1r1w.synth.nz.mem[868] [7];
  assign _09100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [7] : \MSYNC_1r1w.synth.nz.mem[870] [7];
  assign _09101_ = \bapg_rd.w_ptr_r [1] ? _09100_ : _09099_;
  assign _09102_ = \bapg_rd.w_ptr_r [2] ? _09101_ : _09098_;
  assign _09103_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [7] : \MSYNC_1r1w.synth.nz.mem[872] [7];
  assign _09104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [7] : \MSYNC_1r1w.synth.nz.mem[874] [7];
  assign _09105_ = \bapg_rd.w_ptr_r [1] ? _09104_ : _09103_;
  assign _09106_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [7] : \MSYNC_1r1w.synth.nz.mem[876] [7];
  assign _09107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [7] : \MSYNC_1r1w.synth.nz.mem[878] [7];
  assign _09108_ = \bapg_rd.w_ptr_r [1] ? _09107_ : _09106_;
  assign _09109_ = \bapg_rd.w_ptr_r [2] ? _09108_ : _09105_;
  assign _09110_ = \bapg_rd.w_ptr_r [3] ? _09109_ : _09102_;
  assign _09111_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [7] : \MSYNC_1r1w.synth.nz.mem[880] [7];
  assign _09112_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [7] : \MSYNC_1r1w.synth.nz.mem[882] [7];
  assign _09113_ = \bapg_rd.w_ptr_r [1] ? _09112_ : _09111_;
  assign _09114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [7] : \MSYNC_1r1w.synth.nz.mem[884] [7];
  assign _09115_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [7] : \MSYNC_1r1w.synth.nz.mem[886] [7];
  assign _09116_ = \bapg_rd.w_ptr_r [1] ? _09115_ : _09114_;
  assign _09117_ = \bapg_rd.w_ptr_r [2] ? _09116_ : _09113_;
  assign _09118_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [7] : \MSYNC_1r1w.synth.nz.mem[888] [7];
  assign _09119_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [7] : \MSYNC_1r1w.synth.nz.mem[890] [7];
  assign _09120_ = \bapg_rd.w_ptr_r [1] ? _09119_ : _09118_;
  assign _09121_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [7] : \MSYNC_1r1w.synth.nz.mem[892] [7];
  assign _09122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [7] : \MSYNC_1r1w.synth.nz.mem[894] [7];
  assign _09123_ = \bapg_rd.w_ptr_r [1] ? _09122_ : _09121_;
  assign _09124_ = \bapg_rd.w_ptr_r [2] ? _09123_ : _09120_;
  assign _09125_ = \bapg_rd.w_ptr_r [3] ? _09124_ : _09117_;
  assign _09126_ = \bapg_rd.w_ptr_r [4] ? _09125_ : _09110_;
  assign _09127_ = \bapg_rd.w_ptr_r [5] ? _09126_ : _09095_;
  assign _09128_ = \bapg_rd.w_ptr_r [6] ? _09127_ : _09064_;
  assign _09129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [7] : \MSYNC_1r1w.synth.nz.mem[896] [7];
  assign _09130_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [7] : \MSYNC_1r1w.synth.nz.mem[898] [7];
  assign _09131_ = \bapg_rd.w_ptr_r [1] ? _09130_ : _09129_;
  assign _09132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [7] : \MSYNC_1r1w.synth.nz.mem[900] [7];
  assign _09133_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [7] : \MSYNC_1r1w.synth.nz.mem[902] [7];
  assign _09134_ = \bapg_rd.w_ptr_r [1] ? _09133_ : _09132_;
  assign _09135_ = \bapg_rd.w_ptr_r [2] ? _09134_ : _09131_;
  assign _09136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [7] : \MSYNC_1r1w.synth.nz.mem[904] [7];
  assign _09137_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [7] : \MSYNC_1r1w.synth.nz.mem[906] [7];
  assign _09138_ = \bapg_rd.w_ptr_r [1] ? _09137_ : _09136_;
  assign _09139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [7] : \MSYNC_1r1w.synth.nz.mem[908] [7];
  assign _09140_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [7] : \MSYNC_1r1w.synth.nz.mem[910] [7];
  assign _09141_ = \bapg_rd.w_ptr_r [1] ? _09140_ : _09139_;
  assign _09142_ = \bapg_rd.w_ptr_r [2] ? _09141_ : _09138_;
  assign _09143_ = \bapg_rd.w_ptr_r [3] ? _09142_ : _09135_;
  assign _09144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [7] : \MSYNC_1r1w.synth.nz.mem[912] [7];
  assign _09145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [7] : \MSYNC_1r1w.synth.nz.mem[914] [7];
  assign _09146_ = \bapg_rd.w_ptr_r [1] ? _09145_ : _09144_;
  assign _09147_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [7] : \MSYNC_1r1w.synth.nz.mem[916] [7];
  assign _09148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [7] : \MSYNC_1r1w.synth.nz.mem[918] [7];
  assign _09149_ = \bapg_rd.w_ptr_r [1] ? _09148_ : _09147_;
  assign _09150_ = \bapg_rd.w_ptr_r [2] ? _09149_ : _09146_;
  assign _09151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [7] : \MSYNC_1r1w.synth.nz.mem[920] [7];
  assign _09152_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [7] : \MSYNC_1r1w.synth.nz.mem[922] [7];
  assign _09153_ = \bapg_rd.w_ptr_r [1] ? _09152_ : _09151_;
  assign _09154_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [7] : \MSYNC_1r1w.synth.nz.mem[924] [7];
  assign _09155_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [7] : \MSYNC_1r1w.synth.nz.mem[926] [7];
  assign _09156_ = \bapg_rd.w_ptr_r [1] ? _09155_ : _09154_;
  assign _09157_ = \bapg_rd.w_ptr_r [2] ? _09156_ : _09153_;
  assign _09158_ = \bapg_rd.w_ptr_r [3] ? _09157_ : _09150_;
  assign _09159_ = \bapg_rd.w_ptr_r [4] ? _09158_ : _09143_;
  assign _09160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [7] : \MSYNC_1r1w.synth.nz.mem[928] [7];
  assign _09161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [7] : \MSYNC_1r1w.synth.nz.mem[930] [7];
  assign _09162_ = \bapg_rd.w_ptr_r [1] ? _09161_ : _09160_;
  assign _09163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [7] : \MSYNC_1r1w.synth.nz.mem[932] [7];
  assign _09164_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [7] : \MSYNC_1r1w.synth.nz.mem[934] [7];
  assign _09165_ = \bapg_rd.w_ptr_r [1] ? _09164_ : _09163_;
  assign _09166_ = \bapg_rd.w_ptr_r [2] ? _09165_ : _09162_;
  assign _09167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [7] : \MSYNC_1r1w.synth.nz.mem[936] [7];
  assign _09168_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [7] : \MSYNC_1r1w.synth.nz.mem[938] [7];
  assign _09169_ = \bapg_rd.w_ptr_r [1] ? _09168_ : _09167_;
  assign _09170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [7] : \MSYNC_1r1w.synth.nz.mem[940] [7];
  assign _09171_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [7] : \MSYNC_1r1w.synth.nz.mem[942] [7];
  assign _09172_ = \bapg_rd.w_ptr_r [1] ? _09171_ : _09170_;
  assign _09173_ = \bapg_rd.w_ptr_r [2] ? _09172_ : _09169_;
  assign _09174_ = \bapg_rd.w_ptr_r [3] ? _09173_ : _09166_;
  assign _09175_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [7] : \MSYNC_1r1w.synth.nz.mem[944] [7];
  assign _09176_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [7] : \MSYNC_1r1w.synth.nz.mem[946] [7];
  assign _09177_ = \bapg_rd.w_ptr_r [1] ? _09176_ : _09175_;
  assign _09178_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [7] : \MSYNC_1r1w.synth.nz.mem[948] [7];
  assign _09179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [7] : \MSYNC_1r1w.synth.nz.mem[950] [7];
  assign _09180_ = \bapg_rd.w_ptr_r [1] ? _09179_ : _09178_;
  assign _09181_ = \bapg_rd.w_ptr_r [2] ? _09180_ : _09177_;
  assign _09182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [7] : \MSYNC_1r1w.synth.nz.mem[952] [7];
  assign _09183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [7] : \MSYNC_1r1w.synth.nz.mem[954] [7];
  assign _09184_ = \bapg_rd.w_ptr_r [1] ? _09183_ : _09182_;
  assign _09185_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [7] : \MSYNC_1r1w.synth.nz.mem[956] [7];
  assign _09186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [7] : \MSYNC_1r1w.synth.nz.mem[958] [7];
  assign _09187_ = \bapg_rd.w_ptr_r [1] ? _09186_ : _09185_;
  assign _09188_ = \bapg_rd.w_ptr_r [2] ? _09187_ : _09184_;
  assign _09189_ = \bapg_rd.w_ptr_r [3] ? _09188_ : _09181_;
  assign _09190_ = \bapg_rd.w_ptr_r [4] ? _09189_ : _09174_;
  assign _09191_ = \bapg_rd.w_ptr_r [5] ? _09190_ : _09159_;
  assign _09192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [7] : \MSYNC_1r1w.synth.nz.mem[960] [7];
  assign _09193_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [7] : \MSYNC_1r1w.synth.nz.mem[962] [7];
  assign _09194_ = \bapg_rd.w_ptr_r [1] ? _09193_ : _09192_;
  assign _09195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [7] : \MSYNC_1r1w.synth.nz.mem[964] [7];
  assign _09196_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [7] : \MSYNC_1r1w.synth.nz.mem[966] [7];
  assign _09197_ = \bapg_rd.w_ptr_r [1] ? _09196_ : _09195_;
  assign _09198_ = \bapg_rd.w_ptr_r [2] ? _09197_ : _09194_;
  assign _09199_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [7] : \MSYNC_1r1w.synth.nz.mem[968] [7];
  assign _09200_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [7] : \MSYNC_1r1w.synth.nz.mem[970] [7];
  assign _09201_ = \bapg_rd.w_ptr_r [1] ? _09200_ : _09199_;
  assign _09202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [7] : \MSYNC_1r1w.synth.nz.mem[972] [7];
  assign _09203_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [7] : \MSYNC_1r1w.synth.nz.mem[974] [7];
  assign _09204_ = \bapg_rd.w_ptr_r [1] ? _09203_ : _09202_;
  assign _09205_ = \bapg_rd.w_ptr_r [2] ? _09204_ : _09201_;
  assign _09206_ = \bapg_rd.w_ptr_r [3] ? _09205_ : _09198_;
  assign _09207_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [7] : \MSYNC_1r1w.synth.nz.mem[976] [7];
  assign _09208_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [7] : \MSYNC_1r1w.synth.nz.mem[978] [7];
  assign _09209_ = \bapg_rd.w_ptr_r [1] ? _09208_ : _09207_;
  assign _09210_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [7] : \MSYNC_1r1w.synth.nz.mem[980] [7];
  assign _09211_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [7] : \MSYNC_1r1w.synth.nz.mem[982] [7];
  assign _09212_ = \bapg_rd.w_ptr_r [1] ? _09211_ : _09210_;
  assign _09213_ = \bapg_rd.w_ptr_r [2] ? _09212_ : _09209_;
  assign _09214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [7] : \MSYNC_1r1w.synth.nz.mem[984] [7];
  assign _09215_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [7] : \MSYNC_1r1w.synth.nz.mem[986] [7];
  assign _09216_ = \bapg_rd.w_ptr_r [1] ? _09215_ : _09214_;
  assign _09217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [7] : \MSYNC_1r1w.synth.nz.mem[988] [7];
  assign _09218_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [7] : \MSYNC_1r1w.synth.nz.mem[990] [7];
  assign _09219_ = \bapg_rd.w_ptr_r [1] ? _09218_ : _09217_;
  assign _09220_ = \bapg_rd.w_ptr_r [2] ? _09219_ : _09216_;
  assign _09221_ = \bapg_rd.w_ptr_r [3] ? _09220_ : _09213_;
  assign _09222_ = \bapg_rd.w_ptr_r [4] ? _09221_ : _09206_;
  assign _09223_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [7] : \MSYNC_1r1w.synth.nz.mem[992] [7];
  assign _09224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [7] : \MSYNC_1r1w.synth.nz.mem[994] [7];
  assign _09225_ = \bapg_rd.w_ptr_r [1] ? _09224_ : _09223_;
  assign _09226_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [7] : \MSYNC_1r1w.synth.nz.mem[996] [7];
  assign _09227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [7] : \MSYNC_1r1w.synth.nz.mem[998] [7];
  assign _09228_ = \bapg_rd.w_ptr_r [1] ? _09227_ : _09226_;
  assign _09229_ = \bapg_rd.w_ptr_r [2] ? _09228_ : _09225_;
  assign _09230_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [7] : \MSYNC_1r1w.synth.nz.mem[1000] [7];
  assign _09231_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [7] : \MSYNC_1r1w.synth.nz.mem[1002] [7];
  assign _09232_ = \bapg_rd.w_ptr_r [1] ? _09231_ : _09230_;
  assign _09233_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [7] : \MSYNC_1r1w.synth.nz.mem[1004] [7];
  assign _09234_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [7] : \MSYNC_1r1w.synth.nz.mem[1006] [7];
  assign _09235_ = \bapg_rd.w_ptr_r [1] ? _09234_ : _09233_;
  assign _09236_ = \bapg_rd.w_ptr_r [2] ? _09235_ : _09232_;
  assign _09237_ = \bapg_rd.w_ptr_r [3] ? _09236_ : _09229_;
  assign _09238_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [7] : \MSYNC_1r1w.synth.nz.mem[1008] [7];
  assign _09239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [7] : \MSYNC_1r1w.synth.nz.mem[1010] [7];
  assign _09240_ = \bapg_rd.w_ptr_r [1] ? _09239_ : _09238_;
  assign _09241_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [7] : \MSYNC_1r1w.synth.nz.mem[1012] [7];
  assign _09242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [7] : \MSYNC_1r1w.synth.nz.mem[1014] [7];
  assign _09243_ = \bapg_rd.w_ptr_r [1] ? _09242_ : _09241_;
  assign _09244_ = \bapg_rd.w_ptr_r [2] ? _09243_ : _09240_;
  assign _09245_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [7] : \MSYNC_1r1w.synth.nz.mem[1016] [7];
  assign _09246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [7] : \MSYNC_1r1w.synth.nz.mem[1018] [7];
  assign _09247_ = \bapg_rd.w_ptr_r [1] ? _09246_ : _09245_;
  assign _09248_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [7] : \MSYNC_1r1w.synth.nz.mem[1020] [7];
  assign _09249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [7] : \MSYNC_1r1w.synth.nz.mem[1022] [7];
  assign _09250_ = \bapg_rd.w_ptr_r [1] ? _09249_ : _09248_;
  assign _09251_ = \bapg_rd.w_ptr_r [2] ? _09250_ : _09247_;
  assign _09252_ = \bapg_rd.w_ptr_r [3] ? _09251_ : _09244_;
  assign _09253_ = \bapg_rd.w_ptr_r [4] ? _09252_ : _09237_;
  assign _09254_ = \bapg_rd.w_ptr_r [5] ? _09253_ : _09222_;
  assign _09255_ = \bapg_rd.w_ptr_r [6] ? _09254_ : _09191_;
  assign _09256_ = \bapg_rd.w_ptr_r [7] ? _09255_ : _09128_;
  assign _09257_ = \bapg_rd.w_ptr_r [8] ? _09256_ : _09001_;
  assign r_data_o[7] = \bapg_rd.w_ptr_r [9] ? _09257_ : _08746_;
  assign _09258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [8] : \MSYNC_1r1w.synth.nz.mem[0] [8];
  assign _09259_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [8] : \MSYNC_1r1w.synth.nz.mem[2] [8];
  assign _09260_ = \bapg_rd.w_ptr_r [1] ? _09259_ : _09258_;
  assign _09261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [8] : \MSYNC_1r1w.synth.nz.mem[4] [8];
  assign _09262_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [8] : \MSYNC_1r1w.synth.nz.mem[6] [8];
  assign _09263_ = \bapg_rd.w_ptr_r [1] ? _09262_ : _09261_;
  assign _09264_ = \bapg_rd.w_ptr_r [2] ? _09263_ : _09260_;
  assign _09265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [8] : \MSYNC_1r1w.synth.nz.mem[8] [8];
  assign _09266_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [8] : \MSYNC_1r1w.synth.nz.mem[10] [8];
  assign _09267_ = \bapg_rd.w_ptr_r [1] ? _09266_ : _09265_;
  assign _09268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [8] : \MSYNC_1r1w.synth.nz.mem[12] [8];
  assign _09269_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [8] : \MSYNC_1r1w.synth.nz.mem[14] [8];
  assign _09270_ = \bapg_rd.w_ptr_r [1] ? _09269_ : _09268_;
  assign _09271_ = \bapg_rd.w_ptr_r [2] ? _09270_ : _09267_;
  assign _09272_ = \bapg_rd.w_ptr_r [3] ? _09271_ : _09264_;
  assign _09273_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [8] : \MSYNC_1r1w.synth.nz.mem[16] [8];
  assign _09274_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [8] : \MSYNC_1r1w.synth.nz.mem[18] [8];
  assign _09275_ = \bapg_rd.w_ptr_r [1] ? _09274_ : _09273_;
  assign _09276_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [8] : \MSYNC_1r1w.synth.nz.mem[20] [8];
  assign _09277_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [8] : \MSYNC_1r1w.synth.nz.mem[22] [8];
  assign _09278_ = \bapg_rd.w_ptr_r [1] ? _09277_ : _09276_;
  assign _09279_ = \bapg_rd.w_ptr_r [2] ? _09278_ : _09275_;
  assign _09280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [8] : \MSYNC_1r1w.synth.nz.mem[24] [8];
  assign _09281_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [8] : \MSYNC_1r1w.synth.nz.mem[26] [8];
  assign _09282_ = \bapg_rd.w_ptr_r [1] ? _09281_ : _09280_;
  assign _09283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [8] : \MSYNC_1r1w.synth.nz.mem[28] [8];
  assign _09284_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [8] : \MSYNC_1r1w.synth.nz.mem[30] [8];
  assign _09285_ = \bapg_rd.w_ptr_r [1] ? _09284_ : _09283_;
  assign _09286_ = \bapg_rd.w_ptr_r [2] ? _09285_ : _09282_;
  assign _09287_ = \bapg_rd.w_ptr_r [3] ? _09286_ : _09279_;
  assign _09288_ = \bapg_rd.w_ptr_r [4] ? _09287_ : _09272_;
  assign _09289_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [8] : \MSYNC_1r1w.synth.nz.mem[32] [8];
  assign _09290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [8] : \MSYNC_1r1w.synth.nz.mem[34] [8];
  assign _09291_ = \bapg_rd.w_ptr_r [1] ? _09290_ : _09289_;
  assign _09292_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [8] : \MSYNC_1r1w.synth.nz.mem[36] [8];
  assign _09293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [8] : \MSYNC_1r1w.synth.nz.mem[38] [8];
  assign _09294_ = \bapg_rd.w_ptr_r [1] ? _09293_ : _09292_;
  assign _09295_ = \bapg_rd.w_ptr_r [2] ? _09294_ : _09291_;
  assign _09296_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [8] : \MSYNC_1r1w.synth.nz.mem[40] [8];
  assign _09297_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [8] : \MSYNC_1r1w.synth.nz.mem[42] [8];
  assign _09298_ = \bapg_rd.w_ptr_r [1] ? _09297_ : _09296_;
  assign _09299_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [8] : \MSYNC_1r1w.synth.nz.mem[44] [8];
  assign _09300_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [8] : \MSYNC_1r1w.synth.nz.mem[46] [8];
  assign _09301_ = \bapg_rd.w_ptr_r [1] ? _09300_ : _09299_;
  assign _09302_ = \bapg_rd.w_ptr_r [2] ? _09301_ : _09298_;
  assign _09303_ = \bapg_rd.w_ptr_r [3] ? _09302_ : _09295_;
  assign _09304_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [8] : \MSYNC_1r1w.synth.nz.mem[48] [8];
  assign _09305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [8] : \MSYNC_1r1w.synth.nz.mem[50] [8];
  assign _09306_ = \bapg_rd.w_ptr_r [1] ? _09305_ : _09304_;
  assign _09307_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [8] : \MSYNC_1r1w.synth.nz.mem[52] [8];
  assign _09308_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [8] : \MSYNC_1r1w.synth.nz.mem[54] [8];
  assign _09309_ = \bapg_rd.w_ptr_r [1] ? _09308_ : _09307_;
  assign _09310_ = \bapg_rd.w_ptr_r [2] ? _09309_ : _09306_;
  assign _09311_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [8] : \MSYNC_1r1w.synth.nz.mem[56] [8];
  assign _09312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [8] : \MSYNC_1r1w.synth.nz.mem[58] [8];
  assign _09313_ = \bapg_rd.w_ptr_r [1] ? _09312_ : _09311_;
  assign _09314_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [8] : \MSYNC_1r1w.synth.nz.mem[60] [8];
  assign _09315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [8] : \MSYNC_1r1w.synth.nz.mem[62] [8];
  assign _09316_ = \bapg_rd.w_ptr_r [1] ? _09315_ : _09314_;
  assign _09317_ = \bapg_rd.w_ptr_r [2] ? _09316_ : _09313_;
  assign _09318_ = \bapg_rd.w_ptr_r [3] ? _09317_ : _09310_;
  assign _09319_ = \bapg_rd.w_ptr_r [4] ? _09318_ : _09303_;
  assign _09320_ = \bapg_rd.w_ptr_r [5] ? _09319_ : _09288_;
  assign _09321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [8] : \MSYNC_1r1w.synth.nz.mem[64] [8];
  assign _09322_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [8] : \MSYNC_1r1w.synth.nz.mem[66] [8];
  assign _09323_ = \bapg_rd.w_ptr_r [1] ? _09322_ : _09321_;
  assign _09324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [8] : \MSYNC_1r1w.synth.nz.mem[68] [8];
  assign _09325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [8] : \MSYNC_1r1w.synth.nz.mem[70] [8];
  assign _09326_ = \bapg_rd.w_ptr_r [1] ? _09325_ : _09324_;
  assign _09327_ = \bapg_rd.w_ptr_r [2] ? _09326_ : _09323_;
  assign _09328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [8] : \MSYNC_1r1w.synth.nz.mem[72] [8];
  assign _09329_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [8] : \MSYNC_1r1w.synth.nz.mem[74] [8];
  assign _09330_ = \bapg_rd.w_ptr_r [1] ? _09329_ : _09328_;
  assign _09331_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [8] : \MSYNC_1r1w.synth.nz.mem[76] [8];
  assign _09332_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [8] : \MSYNC_1r1w.synth.nz.mem[78] [8];
  assign _09333_ = \bapg_rd.w_ptr_r [1] ? _09332_ : _09331_;
  assign _09334_ = \bapg_rd.w_ptr_r [2] ? _09333_ : _09330_;
  assign _09335_ = \bapg_rd.w_ptr_r [3] ? _09334_ : _09327_;
  assign _09336_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [8] : \MSYNC_1r1w.synth.nz.mem[80] [8];
  assign _09337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [8] : \MSYNC_1r1w.synth.nz.mem[82] [8];
  assign _09338_ = \bapg_rd.w_ptr_r [1] ? _09337_ : _09336_;
  assign _09339_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [8] : \MSYNC_1r1w.synth.nz.mem[84] [8];
  assign _09340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [8] : \MSYNC_1r1w.synth.nz.mem[86] [8];
  assign _09341_ = \bapg_rd.w_ptr_r [1] ? _09340_ : _09339_;
  assign _09342_ = \bapg_rd.w_ptr_r [2] ? _09341_ : _09338_;
  assign _09343_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [8] : \MSYNC_1r1w.synth.nz.mem[88] [8];
  assign _09344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [8] : \MSYNC_1r1w.synth.nz.mem[90] [8];
  assign _09345_ = \bapg_rd.w_ptr_r [1] ? _09344_ : _09343_;
  assign _09346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [8] : \MSYNC_1r1w.synth.nz.mem[92] [8];
  assign _09347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [8] : \MSYNC_1r1w.synth.nz.mem[94] [8];
  assign _09348_ = \bapg_rd.w_ptr_r [1] ? _09347_ : _09346_;
  assign _09349_ = \bapg_rd.w_ptr_r [2] ? _09348_ : _09345_;
  assign _09350_ = \bapg_rd.w_ptr_r [3] ? _09349_ : _09342_;
  assign _09351_ = \bapg_rd.w_ptr_r [4] ? _09350_ : _09335_;
  assign _09352_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [8] : \MSYNC_1r1w.synth.nz.mem[96] [8];
  assign _09353_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [8] : \MSYNC_1r1w.synth.nz.mem[98] [8];
  assign _09354_ = \bapg_rd.w_ptr_r [1] ? _09353_ : _09352_;
  assign _09355_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [8] : \MSYNC_1r1w.synth.nz.mem[100] [8];
  assign _09356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [8] : \MSYNC_1r1w.synth.nz.mem[102] [8];
  assign _09357_ = \bapg_rd.w_ptr_r [1] ? _09356_ : _09355_;
  assign _09358_ = \bapg_rd.w_ptr_r [2] ? _09357_ : _09354_;
  assign _09359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [8] : \MSYNC_1r1w.synth.nz.mem[104] [8];
  assign _09360_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [8] : \MSYNC_1r1w.synth.nz.mem[106] [8];
  assign _09361_ = \bapg_rd.w_ptr_r [1] ? _09360_ : _09359_;
  assign _09362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [8] : \MSYNC_1r1w.synth.nz.mem[108] [8];
  assign _09363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [8] : \MSYNC_1r1w.synth.nz.mem[110] [8];
  assign _09364_ = \bapg_rd.w_ptr_r [1] ? _09363_ : _09362_;
  assign _09365_ = \bapg_rd.w_ptr_r [2] ? _09364_ : _09361_;
  assign _09366_ = \bapg_rd.w_ptr_r [3] ? _09365_ : _09358_;
  assign _09367_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [8] : \MSYNC_1r1w.synth.nz.mem[112] [8];
  assign _09368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [8] : \MSYNC_1r1w.synth.nz.mem[114] [8];
  assign _09369_ = \bapg_rd.w_ptr_r [1] ? _09368_ : _09367_;
  assign _09370_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [8] : \MSYNC_1r1w.synth.nz.mem[116] [8];
  assign _09371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [8] : \MSYNC_1r1w.synth.nz.mem[118] [8];
  assign _09372_ = \bapg_rd.w_ptr_r [1] ? _09371_ : _09370_;
  assign _09373_ = \bapg_rd.w_ptr_r [2] ? _09372_ : _09369_;
  assign _09374_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [8] : \MSYNC_1r1w.synth.nz.mem[120] [8];
  assign _09375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [8] : \MSYNC_1r1w.synth.nz.mem[122] [8];
  assign _09376_ = \bapg_rd.w_ptr_r [1] ? _09375_ : _09374_;
  assign _09377_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [8] : \MSYNC_1r1w.synth.nz.mem[124] [8];
  assign _09378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [8] : \MSYNC_1r1w.synth.nz.mem[126] [8];
  assign _09379_ = \bapg_rd.w_ptr_r [1] ? _09378_ : _09377_;
  assign _09380_ = \bapg_rd.w_ptr_r [2] ? _09379_ : _09376_;
  assign _09381_ = \bapg_rd.w_ptr_r [3] ? _09380_ : _09373_;
  assign _09382_ = \bapg_rd.w_ptr_r [4] ? _09381_ : _09366_;
  assign _09383_ = \bapg_rd.w_ptr_r [5] ? _09382_ : _09351_;
  assign _09384_ = \bapg_rd.w_ptr_r [6] ? _09383_ : _09320_;
  assign _09385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [8] : \MSYNC_1r1w.synth.nz.mem[128] [8];
  assign _09386_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [8] : \MSYNC_1r1w.synth.nz.mem[130] [8];
  assign _09387_ = \bapg_rd.w_ptr_r [1] ? _09386_ : _09385_;
  assign _09388_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [8] : \MSYNC_1r1w.synth.nz.mem[132] [8];
  assign _09389_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [8] : \MSYNC_1r1w.synth.nz.mem[134] [8];
  assign _09390_ = \bapg_rd.w_ptr_r [1] ? _09389_ : _09388_;
  assign _09391_ = \bapg_rd.w_ptr_r [2] ? _09390_ : _09387_;
  assign _09392_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [8] : \MSYNC_1r1w.synth.nz.mem[136] [8];
  assign _09393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [8] : \MSYNC_1r1w.synth.nz.mem[138] [8];
  assign _09394_ = \bapg_rd.w_ptr_r [1] ? _09393_ : _09392_;
  assign _09395_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [8] : \MSYNC_1r1w.synth.nz.mem[140] [8];
  assign _09396_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [8] : \MSYNC_1r1w.synth.nz.mem[142] [8];
  assign _09397_ = \bapg_rd.w_ptr_r [1] ? _09396_ : _09395_;
  assign _09398_ = \bapg_rd.w_ptr_r [2] ? _09397_ : _09394_;
  assign _09399_ = \bapg_rd.w_ptr_r [3] ? _09398_ : _09391_;
  assign _09400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [8] : \MSYNC_1r1w.synth.nz.mem[144] [8];
  assign _09401_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [8] : \MSYNC_1r1w.synth.nz.mem[146] [8];
  assign _09402_ = \bapg_rd.w_ptr_r [1] ? _09401_ : _09400_;
  assign _09403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [8] : \MSYNC_1r1w.synth.nz.mem[148] [8];
  assign _09404_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [8] : \MSYNC_1r1w.synth.nz.mem[150] [8];
  assign _09405_ = \bapg_rd.w_ptr_r [1] ? _09404_ : _09403_;
  assign _09406_ = \bapg_rd.w_ptr_r [2] ? _09405_ : _09402_;
  assign _09407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [8] : \MSYNC_1r1w.synth.nz.mem[152] [8];
  assign _09408_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [8] : \MSYNC_1r1w.synth.nz.mem[154] [8];
  assign _09409_ = \bapg_rd.w_ptr_r [1] ? _09408_ : _09407_;
  assign _09410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [8] : \MSYNC_1r1w.synth.nz.mem[156] [8];
  assign _09411_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [8] : \MSYNC_1r1w.synth.nz.mem[158] [8];
  assign _09412_ = \bapg_rd.w_ptr_r [1] ? _09411_ : _09410_;
  assign _09413_ = \bapg_rd.w_ptr_r [2] ? _09412_ : _09409_;
  assign _09414_ = \bapg_rd.w_ptr_r [3] ? _09413_ : _09406_;
  assign _09415_ = \bapg_rd.w_ptr_r [4] ? _09414_ : _09399_;
  assign _09416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [8] : \MSYNC_1r1w.synth.nz.mem[160] [8];
  assign _09417_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [8] : \MSYNC_1r1w.synth.nz.mem[162] [8];
  assign _09418_ = \bapg_rd.w_ptr_r [1] ? _09417_ : _09416_;
  assign _09419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [8] : \MSYNC_1r1w.synth.nz.mem[164] [8];
  assign _09420_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [8] : \MSYNC_1r1w.synth.nz.mem[166] [8];
  assign _09421_ = \bapg_rd.w_ptr_r [1] ? _09420_ : _09419_;
  assign _09422_ = \bapg_rd.w_ptr_r [2] ? _09421_ : _09418_;
  assign _09423_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [8] : \MSYNC_1r1w.synth.nz.mem[168] [8];
  assign _09424_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [8] : \MSYNC_1r1w.synth.nz.mem[170] [8];
  assign _09425_ = \bapg_rd.w_ptr_r [1] ? _09424_ : _09423_;
  assign _09426_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [8] : \MSYNC_1r1w.synth.nz.mem[172] [8];
  assign _09427_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [8] : \MSYNC_1r1w.synth.nz.mem[174] [8];
  assign _09428_ = \bapg_rd.w_ptr_r [1] ? _09427_ : _09426_;
  assign _09429_ = \bapg_rd.w_ptr_r [2] ? _09428_ : _09425_;
  assign _09430_ = \bapg_rd.w_ptr_r [3] ? _09429_ : _09422_;
  assign _09431_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [8] : \MSYNC_1r1w.synth.nz.mem[176] [8];
  assign _09432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [8] : \MSYNC_1r1w.synth.nz.mem[178] [8];
  assign _09433_ = \bapg_rd.w_ptr_r [1] ? _09432_ : _09431_;
  assign _09434_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [8] : \MSYNC_1r1w.synth.nz.mem[180] [8];
  assign _09435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [8] : \MSYNC_1r1w.synth.nz.mem[182] [8];
  assign _09436_ = \bapg_rd.w_ptr_r [1] ? _09435_ : _09434_;
  assign _09437_ = \bapg_rd.w_ptr_r [2] ? _09436_ : _09433_;
  assign _09438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [8] : \MSYNC_1r1w.synth.nz.mem[184] [8];
  assign _09439_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [8] : \MSYNC_1r1w.synth.nz.mem[186] [8];
  assign _09440_ = \bapg_rd.w_ptr_r [1] ? _09439_ : _09438_;
  assign _09441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [8] : \MSYNC_1r1w.synth.nz.mem[188] [8];
  assign _09442_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [8] : \MSYNC_1r1w.synth.nz.mem[190] [8];
  assign _09443_ = \bapg_rd.w_ptr_r [1] ? _09442_ : _09441_;
  assign _09444_ = \bapg_rd.w_ptr_r [2] ? _09443_ : _09440_;
  assign _09445_ = \bapg_rd.w_ptr_r [3] ? _09444_ : _09437_;
  assign _09446_ = \bapg_rd.w_ptr_r [4] ? _09445_ : _09430_;
  assign _09447_ = \bapg_rd.w_ptr_r [5] ? _09446_ : _09415_;
  assign _09448_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [8] : \MSYNC_1r1w.synth.nz.mem[192] [8];
  assign _09449_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [8] : \MSYNC_1r1w.synth.nz.mem[194] [8];
  assign _09450_ = \bapg_rd.w_ptr_r [1] ? _09449_ : _09448_;
  assign _09451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [8] : \MSYNC_1r1w.synth.nz.mem[196] [8];
  assign _09452_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [8] : \MSYNC_1r1w.synth.nz.mem[198] [8];
  assign _09453_ = \bapg_rd.w_ptr_r [1] ? _09452_ : _09451_;
  assign _09454_ = \bapg_rd.w_ptr_r [2] ? _09453_ : _09450_;
  assign _09455_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [8] : \MSYNC_1r1w.synth.nz.mem[200] [8];
  assign _09456_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [8] : \MSYNC_1r1w.synth.nz.mem[202] [8];
  assign _09457_ = \bapg_rd.w_ptr_r [1] ? _09456_ : _09455_;
  assign _09458_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [8] : \MSYNC_1r1w.synth.nz.mem[204] [8];
  assign _09459_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [8] : \MSYNC_1r1w.synth.nz.mem[206] [8];
  assign _09460_ = \bapg_rd.w_ptr_r [1] ? _09459_ : _09458_;
  assign _09461_ = \bapg_rd.w_ptr_r [2] ? _09460_ : _09457_;
  assign _09462_ = \bapg_rd.w_ptr_r [3] ? _09461_ : _09454_;
  assign _09463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [8] : \MSYNC_1r1w.synth.nz.mem[208] [8];
  assign _09464_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [8] : \MSYNC_1r1w.synth.nz.mem[210] [8];
  assign _09465_ = \bapg_rd.w_ptr_r [1] ? _09464_ : _09463_;
  assign _09466_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [8] : \MSYNC_1r1w.synth.nz.mem[212] [8];
  assign _09467_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [8] : \MSYNC_1r1w.synth.nz.mem[214] [8];
  assign _09468_ = \bapg_rd.w_ptr_r [1] ? _09467_ : _09466_;
  assign _09469_ = \bapg_rd.w_ptr_r [2] ? _09468_ : _09465_;
  assign _09470_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [8] : \MSYNC_1r1w.synth.nz.mem[216] [8];
  assign _09471_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [8] : \MSYNC_1r1w.synth.nz.mem[218] [8];
  assign _09472_ = \bapg_rd.w_ptr_r [1] ? _09471_ : _09470_;
  assign _09473_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [8] : \MSYNC_1r1w.synth.nz.mem[220] [8];
  assign _09474_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [8] : \MSYNC_1r1w.synth.nz.mem[222] [8];
  assign _09475_ = \bapg_rd.w_ptr_r [1] ? _09474_ : _09473_;
  assign _09476_ = \bapg_rd.w_ptr_r [2] ? _09475_ : _09472_;
  assign _09477_ = \bapg_rd.w_ptr_r [3] ? _09476_ : _09469_;
  assign _09478_ = \bapg_rd.w_ptr_r [4] ? _09477_ : _09462_;
  assign _09479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [8] : \MSYNC_1r1w.synth.nz.mem[224] [8];
  assign _09480_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [8] : \MSYNC_1r1w.synth.nz.mem[226] [8];
  assign _09481_ = \bapg_rd.w_ptr_r [1] ? _09480_ : _09479_;
  assign _09482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [8] : \MSYNC_1r1w.synth.nz.mem[228] [8];
  assign _09483_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [8] : \MSYNC_1r1w.synth.nz.mem[230] [8];
  assign _09484_ = \bapg_rd.w_ptr_r [1] ? _09483_ : _09482_;
  assign _09485_ = \bapg_rd.w_ptr_r [2] ? _09484_ : _09481_;
  assign _09486_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [8] : \MSYNC_1r1w.synth.nz.mem[232] [8];
  assign _09487_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [8] : \MSYNC_1r1w.synth.nz.mem[234] [8];
  assign _09488_ = \bapg_rd.w_ptr_r [1] ? _09487_ : _09486_;
  assign _09489_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [8] : \MSYNC_1r1w.synth.nz.mem[236] [8];
  assign _09490_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [8] : \MSYNC_1r1w.synth.nz.mem[238] [8];
  assign _09491_ = \bapg_rd.w_ptr_r [1] ? _09490_ : _09489_;
  assign _09492_ = \bapg_rd.w_ptr_r [2] ? _09491_ : _09488_;
  assign _09493_ = \bapg_rd.w_ptr_r [3] ? _09492_ : _09485_;
  assign _09494_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [8] : \MSYNC_1r1w.synth.nz.mem[240] [8];
  assign _09495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [8] : \MSYNC_1r1w.synth.nz.mem[242] [8];
  assign _09496_ = \bapg_rd.w_ptr_r [1] ? _09495_ : _09494_;
  assign _09497_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [8] : \MSYNC_1r1w.synth.nz.mem[244] [8];
  assign _09498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [8] : \MSYNC_1r1w.synth.nz.mem[246] [8];
  assign _09499_ = \bapg_rd.w_ptr_r [1] ? _09498_ : _09497_;
  assign _09500_ = \bapg_rd.w_ptr_r [2] ? _09499_ : _09496_;
  assign _09501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [8] : \MSYNC_1r1w.synth.nz.mem[248] [8];
  assign _09502_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [8] : \MSYNC_1r1w.synth.nz.mem[250] [8];
  assign _09503_ = \bapg_rd.w_ptr_r [1] ? _09502_ : _09501_;
  assign _09504_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [8] : \MSYNC_1r1w.synth.nz.mem[252] [8];
  assign _09505_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [8] : \MSYNC_1r1w.synth.nz.mem[254] [8];
  assign _09506_ = \bapg_rd.w_ptr_r [1] ? _09505_ : _09504_;
  assign _09507_ = \bapg_rd.w_ptr_r [2] ? _09506_ : _09503_;
  assign _09508_ = \bapg_rd.w_ptr_r [3] ? _09507_ : _09500_;
  assign _09509_ = \bapg_rd.w_ptr_r [4] ? _09508_ : _09493_;
  assign _09510_ = \bapg_rd.w_ptr_r [5] ? _09509_ : _09478_;
  assign _09511_ = \bapg_rd.w_ptr_r [6] ? _09510_ : _09447_;
  assign _09512_ = \bapg_rd.w_ptr_r [7] ? _09511_ : _09384_;
  assign _09513_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [8] : \MSYNC_1r1w.synth.nz.mem[256] [8];
  assign _09514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [8] : \MSYNC_1r1w.synth.nz.mem[258] [8];
  assign _09515_ = \bapg_rd.w_ptr_r [1] ? _09514_ : _09513_;
  assign _09516_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [8] : \MSYNC_1r1w.synth.nz.mem[260] [8];
  assign _09517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [8] : \MSYNC_1r1w.synth.nz.mem[262] [8];
  assign _09518_ = \bapg_rd.w_ptr_r [1] ? _09517_ : _09516_;
  assign _09519_ = \bapg_rd.w_ptr_r [2] ? _09518_ : _09515_;
  assign _09520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [8] : \MSYNC_1r1w.synth.nz.mem[264] [8];
  assign _09521_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [8] : \MSYNC_1r1w.synth.nz.mem[266] [8];
  assign _09522_ = \bapg_rd.w_ptr_r [1] ? _09521_ : _09520_;
  assign _09523_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [8] : \MSYNC_1r1w.synth.nz.mem[268] [8];
  assign _09524_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [8] : \MSYNC_1r1w.synth.nz.mem[270] [8];
  assign _09525_ = \bapg_rd.w_ptr_r [1] ? _09524_ : _09523_;
  assign _09526_ = \bapg_rd.w_ptr_r [2] ? _09525_ : _09522_;
  assign _09527_ = \bapg_rd.w_ptr_r [3] ? _09526_ : _09519_;
  assign _09528_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [8] : \MSYNC_1r1w.synth.nz.mem[272] [8];
  assign _09529_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [8] : \MSYNC_1r1w.synth.nz.mem[274] [8];
  assign _09530_ = \bapg_rd.w_ptr_r [1] ? _09529_ : _09528_;
  assign _09531_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [8] : \MSYNC_1r1w.synth.nz.mem[276] [8];
  assign _09532_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [8] : \MSYNC_1r1w.synth.nz.mem[278] [8];
  assign _09533_ = \bapg_rd.w_ptr_r [1] ? _09532_ : _09531_;
  assign _09534_ = \bapg_rd.w_ptr_r [2] ? _09533_ : _09530_;
  assign _09535_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [8] : \MSYNC_1r1w.synth.nz.mem[280] [8];
  assign _09536_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [8] : \MSYNC_1r1w.synth.nz.mem[282] [8];
  assign _09537_ = \bapg_rd.w_ptr_r [1] ? _09536_ : _09535_;
  assign _09538_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [8] : \MSYNC_1r1w.synth.nz.mem[284] [8];
  assign _09539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [8] : \MSYNC_1r1w.synth.nz.mem[286] [8];
  assign _09540_ = \bapg_rd.w_ptr_r [1] ? _09539_ : _09538_;
  assign _09541_ = \bapg_rd.w_ptr_r [2] ? _09540_ : _09537_;
  assign _09542_ = \bapg_rd.w_ptr_r [3] ? _09541_ : _09534_;
  assign _09543_ = \bapg_rd.w_ptr_r [4] ? _09542_ : _09527_;
  assign _09544_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [8] : \MSYNC_1r1w.synth.nz.mem[288] [8];
  assign _09545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [8] : \MSYNC_1r1w.synth.nz.mem[290] [8];
  assign _09546_ = \bapg_rd.w_ptr_r [1] ? _09545_ : _09544_;
  assign _09547_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [8] : \MSYNC_1r1w.synth.nz.mem[292] [8];
  assign _09548_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [8] : \MSYNC_1r1w.synth.nz.mem[294] [8];
  assign _09549_ = \bapg_rd.w_ptr_r [1] ? _09548_ : _09547_;
  assign _09550_ = \bapg_rd.w_ptr_r [2] ? _09549_ : _09546_;
  assign _09551_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [8] : \MSYNC_1r1w.synth.nz.mem[296] [8];
  assign _09552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [8] : \MSYNC_1r1w.synth.nz.mem[298] [8];
  assign _09553_ = \bapg_rd.w_ptr_r [1] ? _09552_ : _09551_;
  assign _09554_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [8] : \MSYNC_1r1w.synth.nz.mem[300] [8];
  assign _09555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [8] : \MSYNC_1r1w.synth.nz.mem[302] [8];
  assign _09556_ = \bapg_rd.w_ptr_r [1] ? _09555_ : _09554_;
  assign _09557_ = \bapg_rd.w_ptr_r [2] ? _09556_ : _09553_;
  assign _09558_ = \bapg_rd.w_ptr_r [3] ? _09557_ : _09550_;
  assign _09559_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [8] : \MSYNC_1r1w.synth.nz.mem[304] [8];
  assign _09560_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [8] : \MSYNC_1r1w.synth.nz.mem[306] [8];
  assign _09561_ = \bapg_rd.w_ptr_r [1] ? _09560_ : _09559_;
  assign _09562_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [8] : \MSYNC_1r1w.synth.nz.mem[308] [8];
  assign _09563_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [8] : \MSYNC_1r1w.synth.nz.mem[310] [8];
  assign _09564_ = \bapg_rd.w_ptr_r [1] ? _09563_ : _09562_;
  assign _09565_ = \bapg_rd.w_ptr_r [2] ? _09564_ : _09561_;
  assign _09566_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [8] : \MSYNC_1r1w.synth.nz.mem[312] [8];
  assign _09567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [8] : \MSYNC_1r1w.synth.nz.mem[314] [8];
  assign _09568_ = \bapg_rd.w_ptr_r [1] ? _09567_ : _09566_;
  assign _09569_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [8] : \MSYNC_1r1w.synth.nz.mem[316] [8];
  assign _09570_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [8] : \MSYNC_1r1w.synth.nz.mem[318] [8];
  assign _09571_ = \bapg_rd.w_ptr_r [1] ? _09570_ : _09569_;
  assign _09572_ = \bapg_rd.w_ptr_r [2] ? _09571_ : _09568_;
  assign _09573_ = \bapg_rd.w_ptr_r [3] ? _09572_ : _09565_;
  assign _09574_ = \bapg_rd.w_ptr_r [4] ? _09573_ : _09558_;
  assign _09575_ = \bapg_rd.w_ptr_r [5] ? _09574_ : _09543_;
  assign _09576_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [8] : \MSYNC_1r1w.synth.nz.mem[320] [8];
  assign _09577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [8] : \MSYNC_1r1w.synth.nz.mem[322] [8];
  assign _09578_ = \bapg_rd.w_ptr_r [1] ? _09577_ : _09576_;
  assign _09579_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [8] : \MSYNC_1r1w.synth.nz.mem[324] [8];
  assign _09580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [8] : \MSYNC_1r1w.synth.nz.mem[326] [8];
  assign _09581_ = \bapg_rd.w_ptr_r [1] ? _09580_ : _09579_;
  assign _09582_ = \bapg_rd.w_ptr_r [2] ? _09581_ : _09578_;
  assign _09583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [8] : \MSYNC_1r1w.synth.nz.mem[328] [8];
  assign _09584_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [8] : \MSYNC_1r1w.synth.nz.mem[330] [8];
  assign _09585_ = \bapg_rd.w_ptr_r [1] ? _09584_ : _09583_;
  assign _09586_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [8] : \MSYNC_1r1w.synth.nz.mem[332] [8];
  assign _09587_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [8] : \MSYNC_1r1w.synth.nz.mem[334] [8];
  assign _09588_ = \bapg_rd.w_ptr_r [1] ? _09587_ : _09586_;
  assign _09589_ = \bapg_rd.w_ptr_r [2] ? _09588_ : _09585_;
  assign _09590_ = \bapg_rd.w_ptr_r [3] ? _09589_ : _09582_;
  assign _09591_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [8] : \MSYNC_1r1w.synth.nz.mem[336] [8];
  assign _09592_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [8] : \MSYNC_1r1w.synth.nz.mem[338] [8];
  assign _09593_ = \bapg_rd.w_ptr_r [1] ? _09592_ : _09591_;
  assign _09594_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [8] : \MSYNC_1r1w.synth.nz.mem[340] [8];
  assign _09595_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [8] : \MSYNC_1r1w.synth.nz.mem[342] [8];
  assign _09596_ = \bapg_rd.w_ptr_r [1] ? _09595_ : _09594_;
  assign _09597_ = \bapg_rd.w_ptr_r [2] ? _09596_ : _09593_;
  assign _09598_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [8] : \MSYNC_1r1w.synth.nz.mem[344] [8];
  assign _09599_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [8] : \MSYNC_1r1w.synth.nz.mem[346] [8];
  assign _09600_ = \bapg_rd.w_ptr_r [1] ? _09599_ : _09598_;
  assign _09601_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [8] : \MSYNC_1r1w.synth.nz.mem[348] [8];
  assign _09602_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [8] : \MSYNC_1r1w.synth.nz.mem[350] [8];
  assign _09603_ = \bapg_rd.w_ptr_r [1] ? _09602_ : _09601_;
  assign _09604_ = \bapg_rd.w_ptr_r [2] ? _09603_ : _09600_;
  assign _09605_ = \bapg_rd.w_ptr_r [3] ? _09604_ : _09597_;
  assign _09606_ = \bapg_rd.w_ptr_r [4] ? _09605_ : _09590_;
  assign _09607_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [8] : \MSYNC_1r1w.synth.nz.mem[352] [8];
  assign _09608_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [8] : \MSYNC_1r1w.synth.nz.mem[354] [8];
  assign _09609_ = \bapg_rd.w_ptr_r [1] ? _09608_ : _09607_;
  assign _09610_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [8] : \MSYNC_1r1w.synth.nz.mem[356] [8];
  assign _09611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [8] : \MSYNC_1r1w.synth.nz.mem[358] [8];
  assign _09612_ = \bapg_rd.w_ptr_r [1] ? _09611_ : _09610_;
  assign _09613_ = \bapg_rd.w_ptr_r [2] ? _09612_ : _09609_;
  assign _09614_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [8] : \MSYNC_1r1w.synth.nz.mem[360] [8];
  assign _09615_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [8] : \MSYNC_1r1w.synth.nz.mem[362] [8];
  assign _09616_ = \bapg_rd.w_ptr_r [1] ? _09615_ : _09614_;
  assign _09617_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [8] : \MSYNC_1r1w.synth.nz.mem[364] [8];
  assign _09618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [8] : \MSYNC_1r1w.synth.nz.mem[366] [8];
  assign _09619_ = \bapg_rd.w_ptr_r [1] ? _09618_ : _09617_;
  assign _09620_ = \bapg_rd.w_ptr_r [2] ? _09619_ : _09616_;
  assign _09621_ = \bapg_rd.w_ptr_r [3] ? _09620_ : _09613_;
  assign _09622_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [8] : \MSYNC_1r1w.synth.nz.mem[368] [8];
  assign _09623_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [8] : \MSYNC_1r1w.synth.nz.mem[370] [8];
  assign _09624_ = \bapg_rd.w_ptr_r [1] ? _09623_ : _09622_;
  assign _09625_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [8] : \MSYNC_1r1w.synth.nz.mem[372] [8];
  assign _09626_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [8] : \MSYNC_1r1w.synth.nz.mem[374] [8];
  assign _09627_ = \bapg_rd.w_ptr_r [1] ? _09626_ : _09625_;
  assign _09628_ = \bapg_rd.w_ptr_r [2] ? _09627_ : _09624_;
  assign _09629_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [8] : \MSYNC_1r1w.synth.nz.mem[376] [8];
  assign _09630_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [8] : \MSYNC_1r1w.synth.nz.mem[378] [8];
  assign _09631_ = \bapg_rd.w_ptr_r [1] ? _09630_ : _09629_;
  assign _09632_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [8] : \MSYNC_1r1w.synth.nz.mem[380] [8];
  assign _09633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [8] : \MSYNC_1r1w.synth.nz.mem[382] [8];
  assign _09634_ = \bapg_rd.w_ptr_r [1] ? _09633_ : _09632_;
  assign _09635_ = \bapg_rd.w_ptr_r [2] ? _09634_ : _09631_;
  assign _09636_ = \bapg_rd.w_ptr_r [3] ? _09635_ : _09628_;
  assign _09637_ = \bapg_rd.w_ptr_r [4] ? _09636_ : _09621_;
  assign _09638_ = \bapg_rd.w_ptr_r [5] ? _09637_ : _09606_;
  assign _09639_ = \bapg_rd.w_ptr_r [6] ? _09638_ : _09575_;
  assign _09640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [8] : \MSYNC_1r1w.synth.nz.mem[384] [8];
  assign _09641_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [8] : \MSYNC_1r1w.synth.nz.mem[386] [8];
  assign _09642_ = \bapg_rd.w_ptr_r [1] ? _09641_ : _09640_;
  assign _09643_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [8] : \MSYNC_1r1w.synth.nz.mem[388] [8];
  assign _09644_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [8] : \MSYNC_1r1w.synth.nz.mem[390] [8];
  assign _09645_ = \bapg_rd.w_ptr_r [1] ? _09644_ : _09643_;
  assign _09646_ = \bapg_rd.w_ptr_r [2] ? _09645_ : _09642_;
  assign _09647_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [8] : \MSYNC_1r1w.synth.nz.mem[392] [8];
  assign _09648_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [8] : \MSYNC_1r1w.synth.nz.mem[394] [8];
  assign _09649_ = \bapg_rd.w_ptr_r [1] ? _09648_ : _09647_;
  assign _09650_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [8] : \MSYNC_1r1w.synth.nz.mem[396] [8];
  assign _09651_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [8] : \MSYNC_1r1w.synth.nz.mem[398] [8];
  assign _09652_ = \bapg_rd.w_ptr_r [1] ? _09651_ : _09650_;
  assign _09653_ = \bapg_rd.w_ptr_r [2] ? _09652_ : _09649_;
  assign _09654_ = \bapg_rd.w_ptr_r [3] ? _09653_ : _09646_;
  assign _09655_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [8] : \MSYNC_1r1w.synth.nz.mem[400] [8];
  assign _09656_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [8] : \MSYNC_1r1w.synth.nz.mem[402] [8];
  assign _09657_ = \bapg_rd.w_ptr_r [1] ? _09656_ : _09655_;
  assign _09658_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [8] : \MSYNC_1r1w.synth.nz.mem[404] [8];
  assign _09659_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [8] : \MSYNC_1r1w.synth.nz.mem[406] [8];
  assign _09660_ = \bapg_rd.w_ptr_r [1] ? _09659_ : _09658_;
  assign _09661_ = \bapg_rd.w_ptr_r [2] ? _09660_ : _09657_;
  assign _09662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [8] : \MSYNC_1r1w.synth.nz.mem[408] [8];
  assign _09663_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [8] : \MSYNC_1r1w.synth.nz.mem[410] [8];
  assign _09664_ = \bapg_rd.w_ptr_r [1] ? _09663_ : _09662_;
  assign _09665_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [8] : \MSYNC_1r1w.synth.nz.mem[412] [8];
  assign _09666_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [8] : \MSYNC_1r1w.synth.nz.mem[414] [8];
  assign _09667_ = \bapg_rd.w_ptr_r [1] ? _09666_ : _09665_;
  assign _09668_ = \bapg_rd.w_ptr_r [2] ? _09667_ : _09664_;
  assign _09669_ = \bapg_rd.w_ptr_r [3] ? _09668_ : _09661_;
  assign _09670_ = \bapg_rd.w_ptr_r [4] ? _09669_ : _09654_;
  assign _09671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [8] : \MSYNC_1r1w.synth.nz.mem[416] [8];
  assign _09672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [8] : \MSYNC_1r1w.synth.nz.mem[418] [8];
  assign _09673_ = \bapg_rd.w_ptr_r [1] ? _09672_ : _09671_;
  assign _09674_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [8] : \MSYNC_1r1w.synth.nz.mem[420] [8];
  assign _09675_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [8] : \MSYNC_1r1w.synth.nz.mem[422] [8];
  assign _09676_ = \bapg_rd.w_ptr_r [1] ? _09675_ : _09674_;
  assign _09677_ = \bapg_rd.w_ptr_r [2] ? _09676_ : _09673_;
  assign _09678_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [8] : \MSYNC_1r1w.synth.nz.mem[424] [8];
  assign _09679_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [8] : \MSYNC_1r1w.synth.nz.mem[426] [8];
  assign _09680_ = \bapg_rd.w_ptr_r [1] ? _09679_ : _09678_;
  assign _09681_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [8] : \MSYNC_1r1w.synth.nz.mem[428] [8];
  assign _09682_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [8] : \MSYNC_1r1w.synth.nz.mem[430] [8];
  assign _09683_ = \bapg_rd.w_ptr_r [1] ? _09682_ : _09681_;
  assign _09684_ = \bapg_rd.w_ptr_r [2] ? _09683_ : _09680_;
  assign _09685_ = \bapg_rd.w_ptr_r [3] ? _09684_ : _09677_;
  assign _09686_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [8] : \MSYNC_1r1w.synth.nz.mem[432] [8];
  assign _09687_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [8] : \MSYNC_1r1w.synth.nz.mem[434] [8];
  assign _09688_ = \bapg_rd.w_ptr_r [1] ? _09687_ : _09686_;
  assign _09689_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [8] : \MSYNC_1r1w.synth.nz.mem[436] [8];
  assign _09690_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [8] : \MSYNC_1r1w.synth.nz.mem[438] [8];
  assign _09691_ = \bapg_rd.w_ptr_r [1] ? _09690_ : _09689_;
  assign _09692_ = \bapg_rd.w_ptr_r [2] ? _09691_ : _09688_;
  assign _09693_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [8] : \MSYNC_1r1w.synth.nz.mem[440] [8];
  assign _09694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [8] : \MSYNC_1r1w.synth.nz.mem[442] [8];
  assign _09695_ = \bapg_rd.w_ptr_r [1] ? _09694_ : _09693_;
  assign _09696_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [8] : \MSYNC_1r1w.synth.nz.mem[444] [8];
  assign _09697_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [8] : \MSYNC_1r1w.synth.nz.mem[446] [8];
  assign _09698_ = \bapg_rd.w_ptr_r [1] ? _09697_ : _09696_;
  assign _09699_ = \bapg_rd.w_ptr_r [2] ? _09698_ : _09695_;
  assign _09700_ = \bapg_rd.w_ptr_r [3] ? _09699_ : _09692_;
  assign _09701_ = \bapg_rd.w_ptr_r [4] ? _09700_ : _09685_;
  assign _09702_ = \bapg_rd.w_ptr_r [5] ? _09701_ : _09670_;
  assign _09703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [8] : \MSYNC_1r1w.synth.nz.mem[448] [8];
  assign _09704_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [8] : \MSYNC_1r1w.synth.nz.mem[450] [8];
  assign _09705_ = \bapg_rd.w_ptr_r [1] ? _09704_ : _09703_;
  assign _09706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [8] : \MSYNC_1r1w.synth.nz.mem[452] [8];
  assign _09707_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [8] : \MSYNC_1r1w.synth.nz.mem[454] [8];
  assign _09708_ = \bapg_rd.w_ptr_r [1] ? _09707_ : _09706_;
  assign _09709_ = \bapg_rd.w_ptr_r [2] ? _09708_ : _09705_;
  assign _09710_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [8] : \MSYNC_1r1w.synth.nz.mem[456] [8];
  assign _09711_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [8] : \MSYNC_1r1w.synth.nz.mem[458] [8];
  assign _09712_ = \bapg_rd.w_ptr_r [1] ? _09711_ : _09710_;
  assign _09713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [8] : \MSYNC_1r1w.synth.nz.mem[460] [8];
  assign _09714_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [8] : \MSYNC_1r1w.synth.nz.mem[462] [8];
  assign _09715_ = \bapg_rd.w_ptr_r [1] ? _09714_ : _09713_;
  assign _09716_ = \bapg_rd.w_ptr_r [2] ? _09715_ : _09712_;
  assign _09717_ = \bapg_rd.w_ptr_r [3] ? _09716_ : _09709_;
  assign _09718_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [8] : \MSYNC_1r1w.synth.nz.mem[464] [8];
  assign _09719_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [8] : \MSYNC_1r1w.synth.nz.mem[466] [8];
  assign _09720_ = \bapg_rd.w_ptr_r [1] ? _09719_ : _09718_;
  assign _09721_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [8] : \MSYNC_1r1w.synth.nz.mem[468] [8];
  assign _09722_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [8] : \MSYNC_1r1w.synth.nz.mem[470] [8];
  assign _09723_ = \bapg_rd.w_ptr_r [1] ? _09722_ : _09721_;
  assign _09724_ = \bapg_rd.w_ptr_r [2] ? _09723_ : _09720_;
  assign _09725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [8] : \MSYNC_1r1w.synth.nz.mem[472] [8];
  assign _09726_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [8] : \MSYNC_1r1w.synth.nz.mem[474] [8];
  assign _09727_ = \bapg_rd.w_ptr_r [1] ? _09726_ : _09725_;
  assign _09728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [8] : \MSYNC_1r1w.synth.nz.mem[476] [8];
  assign _09729_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [8] : \MSYNC_1r1w.synth.nz.mem[478] [8];
  assign _09730_ = \bapg_rd.w_ptr_r [1] ? _09729_ : _09728_;
  assign _09731_ = \bapg_rd.w_ptr_r [2] ? _09730_ : _09727_;
  assign _09732_ = \bapg_rd.w_ptr_r [3] ? _09731_ : _09724_;
  assign _09733_ = \bapg_rd.w_ptr_r [4] ? _09732_ : _09717_;
  assign _09734_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [8] : \MSYNC_1r1w.synth.nz.mem[480] [8];
  assign _09735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [8] : \MSYNC_1r1w.synth.nz.mem[482] [8];
  assign _09736_ = \bapg_rd.w_ptr_r [1] ? _09735_ : _09734_;
  assign _09737_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [8] : \MSYNC_1r1w.synth.nz.mem[484] [8];
  assign _09738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [8] : \MSYNC_1r1w.synth.nz.mem[486] [8];
  assign _09739_ = \bapg_rd.w_ptr_r [1] ? _09738_ : _09737_;
  assign _09740_ = \bapg_rd.w_ptr_r [2] ? _09739_ : _09736_;
  assign _09741_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [8] : \MSYNC_1r1w.synth.nz.mem[488] [8];
  assign _09742_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [8] : \MSYNC_1r1w.synth.nz.mem[490] [8];
  assign _09743_ = \bapg_rd.w_ptr_r [1] ? _09742_ : _09741_;
  assign _09744_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [8] : \MSYNC_1r1w.synth.nz.mem[492] [8];
  assign _09745_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [8] : \MSYNC_1r1w.synth.nz.mem[494] [8];
  assign _09746_ = \bapg_rd.w_ptr_r [1] ? _09745_ : _09744_;
  assign _09747_ = \bapg_rd.w_ptr_r [2] ? _09746_ : _09743_;
  assign _09748_ = \bapg_rd.w_ptr_r [3] ? _09747_ : _09740_;
  assign _09749_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [8] : \MSYNC_1r1w.synth.nz.mem[496] [8];
  assign _09750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [8] : \MSYNC_1r1w.synth.nz.mem[498] [8];
  assign _09751_ = \bapg_rd.w_ptr_r [1] ? _09750_ : _09749_;
  assign _09752_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [8] : \MSYNC_1r1w.synth.nz.mem[500] [8];
  assign _09753_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [8] : \MSYNC_1r1w.synth.nz.mem[502] [8];
  assign _09754_ = \bapg_rd.w_ptr_r [1] ? _09753_ : _09752_;
  assign _09755_ = \bapg_rd.w_ptr_r [2] ? _09754_ : _09751_;
  assign _09756_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [8] : \MSYNC_1r1w.synth.nz.mem[504] [8];
  assign _09757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [8] : \MSYNC_1r1w.synth.nz.mem[506] [8];
  assign _09758_ = \bapg_rd.w_ptr_r [1] ? _09757_ : _09756_;
  assign _09759_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [8] : \MSYNC_1r1w.synth.nz.mem[508] [8];
  assign _09760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [8] : \MSYNC_1r1w.synth.nz.mem[510] [8];
  assign _09761_ = \bapg_rd.w_ptr_r [1] ? _09760_ : _09759_;
  assign _09762_ = \bapg_rd.w_ptr_r [2] ? _09761_ : _09758_;
  assign _09763_ = \bapg_rd.w_ptr_r [3] ? _09762_ : _09755_;
  assign _09764_ = \bapg_rd.w_ptr_r [4] ? _09763_ : _09748_;
  assign _09765_ = \bapg_rd.w_ptr_r [5] ? _09764_ : _09733_;
  assign _09766_ = \bapg_rd.w_ptr_r [6] ? _09765_ : _09702_;
  assign _09767_ = \bapg_rd.w_ptr_r [7] ? _09766_ : _09639_;
  assign _09768_ = \bapg_rd.w_ptr_r [8] ? _09767_ : _09512_;
  assign _09769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [8] : \MSYNC_1r1w.synth.nz.mem[512] [8];
  assign _09770_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [8] : \MSYNC_1r1w.synth.nz.mem[514] [8];
  assign _09771_ = \bapg_rd.w_ptr_r [1] ? _09770_ : _09769_;
  assign _09772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [8] : \MSYNC_1r1w.synth.nz.mem[516] [8];
  assign _09773_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [8] : \MSYNC_1r1w.synth.nz.mem[518] [8];
  assign _09774_ = \bapg_rd.w_ptr_r [1] ? _09773_ : _09772_;
  assign _09775_ = \bapg_rd.w_ptr_r [2] ? _09774_ : _09771_;
  assign _09776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [8] : \MSYNC_1r1w.synth.nz.mem[520] [8];
  assign _09777_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [8] : \MSYNC_1r1w.synth.nz.mem[522] [8];
  assign _09778_ = \bapg_rd.w_ptr_r [1] ? _09777_ : _09776_;
  assign _09779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [8] : \MSYNC_1r1w.synth.nz.mem[524] [8];
  assign _09780_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [8] : \MSYNC_1r1w.synth.nz.mem[526] [8];
  assign _09781_ = \bapg_rd.w_ptr_r [1] ? _09780_ : _09779_;
  assign _09782_ = \bapg_rd.w_ptr_r [2] ? _09781_ : _09778_;
  assign _09783_ = \bapg_rd.w_ptr_r [3] ? _09782_ : _09775_;
  assign _09784_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [8] : \MSYNC_1r1w.synth.nz.mem[528] [8];
  assign _09785_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [8] : \MSYNC_1r1w.synth.nz.mem[530] [8];
  assign _09786_ = \bapg_rd.w_ptr_r [1] ? _09785_ : _09784_;
  assign _09787_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [8] : \MSYNC_1r1w.synth.nz.mem[532] [8];
  assign _09788_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [8] : \MSYNC_1r1w.synth.nz.mem[534] [8];
  assign _09789_ = \bapg_rd.w_ptr_r [1] ? _09788_ : _09787_;
  assign _09790_ = \bapg_rd.w_ptr_r [2] ? _09789_ : _09786_;
  assign _09791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [8] : \MSYNC_1r1w.synth.nz.mem[536] [8];
  assign _09792_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [8] : \MSYNC_1r1w.synth.nz.mem[538] [8];
  assign _09793_ = \bapg_rd.w_ptr_r [1] ? _09792_ : _09791_;
  assign _09794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [8] : \MSYNC_1r1w.synth.nz.mem[540] [8];
  assign _09795_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [8] : \MSYNC_1r1w.synth.nz.mem[542] [8];
  assign _09796_ = \bapg_rd.w_ptr_r [1] ? _09795_ : _09794_;
  assign _09797_ = \bapg_rd.w_ptr_r [2] ? _09796_ : _09793_;
  assign _09798_ = \bapg_rd.w_ptr_r [3] ? _09797_ : _09790_;
  assign _09799_ = \bapg_rd.w_ptr_r [4] ? _09798_ : _09783_;
  assign _09800_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [8] : \MSYNC_1r1w.synth.nz.mem[544] [8];
  assign _09801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [8] : \MSYNC_1r1w.synth.nz.mem[546] [8];
  assign _09802_ = \bapg_rd.w_ptr_r [1] ? _09801_ : _09800_;
  assign _09803_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [8] : \MSYNC_1r1w.synth.nz.mem[548] [8];
  assign _09804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [8] : \MSYNC_1r1w.synth.nz.mem[550] [8];
  assign _09805_ = \bapg_rd.w_ptr_r [1] ? _09804_ : _09803_;
  assign _09806_ = \bapg_rd.w_ptr_r [2] ? _09805_ : _09802_;
  assign _09807_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [8] : \MSYNC_1r1w.synth.nz.mem[552] [8];
  assign _09808_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [8] : \MSYNC_1r1w.synth.nz.mem[554] [8];
  assign _09809_ = \bapg_rd.w_ptr_r [1] ? _09808_ : _09807_;
  assign _09810_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [8] : \MSYNC_1r1w.synth.nz.mem[556] [8];
  assign _09811_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [8] : \MSYNC_1r1w.synth.nz.mem[558] [8];
  assign _09812_ = \bapg_rd.w_ptr_r [1] ? _09811_ : _09810_;
  assign _09813_ = \bapg_rd.w_ptr_r [2] ? _09812_ : _09809_;
  assign _09814_ = \bapg_rd.w_ptr_r [3] ? _09813_ : _09806_;
  assign _09815_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [8] : \MSYNC_1r1w.synth.nz.mem[560] [8];
  assign _09816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [8] : \MSYNC_1r1w.synth.nz.mem[562] [8];
  assign _09817_ = \bapg_rd.w_ptr_r [1] ? _09816_ : _09815_;
  assign _09818_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [8] : \MSYNC_1r1w.synth.nz.mem[564] [8];
  assign _09819_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [8] : \MSYNC_1r1w.synth.nz.mem[566] [8];
  assign _09820_ = \bapg_rd.w_ptr_r [1] ? _09819_ : _09818_;
  assign _09821_ = \bapg_rd.w_ptr_r [2] ? _09820_ : _09817_;
  assign _09822_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [8] : \MSYNC_1r1w.synth.nz.mem[568] [8];
  assign _09823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [8] : \MSYNC_1r1w.synth.nz.mem[570] [8];
  assign _09824_ = \bapg_rd.w_ptr_r [1] ? _09823_ : _09822_;
  assign _09825_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [8] : \MSYNC_1r1w.synth.nz.mem[572] [8];
  assign _09826_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [8] : \MSYNC_1r1w.synth.nz.mem[574] [8];
  assign _09827_ = \bapg_rd.w_ptr_r [1] ? _09826_ : _09825_;
  assign _09828_ = \bapg_rd.w_ptr_r [2] ? _09827_ : _09824_;
  assign _09829_ = \bapg_rd.w_ptr_r [3] ? _09828_ : _09821_;
  assign _09830_ = \bapg_rd.w_ptr_r [4] ? _09829_ : _09814_;
  assign _09831_ = \bapg_rd.w_ptr_r [5] ? _09830_ : _09799_;
  assign _09832_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [8] : \MSYNC_1r1w.synth.nz.mem[576] [8];
  assign _09833_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [8] : \MSYNC_1r1w.synth.nz.mem[578] [8];
  assign _09834_ = \bapg_rd.w_ptr_r [1] ? _09833_ : _09832_;
  assign _09835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [8] : \MSYNC_1r1w.synth.nz.mem[580] [8];
  assign _09836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [8] : \MSYNC_1r1w.synth.nz.mem[582] [8];
  assign _09837_ = \bapg_rd.w_ptr_r [1] ? _09836_ : _09835_;
  assign _09838_ = \bapg_rd.w_ptr_r [2] ? _09837_ : _09834_;
  assign _09839_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [8] : \MSYNC_1r1w.synth.nz.mem[584] [8];
  assign _09840_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [8] : \MSYNC_1r1w.synth.nz.mem[586] [8];
  assign _09841_ = \bapg_rd.w_ptr_r [1] ? _09840_ : _09839_;
  assign _09842_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [8] : \MSYNC_1r1w.synth.nz.mem[588] [8];
  assign _09843_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [8] : \MSYNC_1r1w.synth.nz.mem[590] [8];
  assign _09844_ = \bapg_rd.w_ptr_r [1] ? _09843_ : _09842_;
  assign _09845_ = \bapg_rd.w_ptr_r [2] ? _09844_ : _09841_;
  assign _09846_ = \bapg_rd.w_ptr_r [3] ? _09845_ : _09838_;
  assign _09847_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [8] : \MSYNC_1r1w.synth.nz.mem[592] [8];
  assign _09848_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [8] : \MSYNC_1r1w.synth.nz.mem[594] [8];
  assign _09849_ = \bapg_rd.w_ptr_r [1] ? _09848_ : _09847_;
  assign _09850_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [8] : \MSYNC_1r1w.synth.nz.mem[596] [8];
  assign _09851_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [8] : \MSYNC_1r1w.synth.nz.mem[598] [8];
  assign _09852_ = \bapg_rd.w_ptr_r [1] ? _09851_ : _09850_;
  assign _09853_ = \bapg_rd.w_ptr_r [2] ? _09852_ : _09849_;
  assign _09854_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [8] : \MSYNC_1r1w.synth.nz.mem[600] [8];
  assign _09855_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [8] : \MSYNC_1r1w.synth.nz.mem[602] [8];
  assign _09856_ = \bapg_rd.w_ptr_r [1] ? _09855_ : _09854_;
  assign _09857_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [8] : \MSYNC_1r1w.synth.nz.mem[604] [8];
  assign _09858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [8] : \MSYNC_1r1w.synth.nz.mem[606] [8];
  assign _09859_ = \bapg_rd.w_ptr_r [1] ? _09858_ : _09857_;
  assign _09860_ = \bapg_rd.w_ptr_r [2] ? _09859_ : _09856_;
  assign _09861_ = \bapg_rd.w_ptr_r [3] ? _09860_ : _09853_;
  assign _09862_ = \bapg_rd.w_ptr_r [4] ? _09861_ : _09846_;
  assign _09863_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [8] : \MSYNC_1r1w.synth.nz.mem[608] [8];
  assign _09864_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [8] : \MSYNC_1r1w.synth.nz.mem[610] [8];
  assign _09865_ = \bapg_rd.w_ptr_r [1] ? _09864_ : _09863_;
  assign _09866_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [8] : \MSYNC_1r1w.synth.nz.mem[612] [8];
  assign _09867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [8] : \MSYNC_1r1w.synth.nz.mem[614] [8];
  assign _09868_ = \bapg_rd.w_ptr_r [1] ? _09867_ : _09866_;
  assign _09869_ = \bapg_rd.w_ptr_r [2] ? _09868_ : _09865_;
  assign _09870_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [8] : \MSYNC_1r1w.synth.nz.mem[616] [8];
  assign _09871_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [8] : \MSYNC_1r1w.synth.nz.mem[618] [8];
  assign _09872_ = \bapg_rd.w_ptr_r [1] ? _09871_ : _09870_;
  assign _09873_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [8] : \MSYNC_1r1w.synth.nz.mem[620] [8];
  assign _09874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [8] : \MSYNC_1r1w.synth.nz.mem[622] [8];
  assign _09875_ = \bapg_rd.w_ptr_r [1] ? _09874_ : _09873_;
  assign _09876_ = \bapg_rd.w_ptr_r [2] ? _09875_ : _09872_;
  assign _09877_ = \bapg_rd.w_ptr_r [3] ? _09876_ : _09869_;
  assign _09878_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [8] : \MSYNC_1r1w.synth.nz.mem[624] [8];
  assign _09879_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [8] : \MSYNC_1r1w.synth.nz.mem[626] [8];
  assign _09880_ = \bapg_rd.w_ptr_r [1] ? _09879_ : _09878_;
  assign _09881_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [8] : \MSYNC_1r1w.synth.nz.mem[628] [8];
  assign _09882_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [8] : \MSYNC_1r1w.synth.nz.mem[630] [8];
  assign _09883_ = \bapg_rd.w_ptr_r [1] ? _09882_ : _09881_;
  assign _09884_ = \bapg_rd.w_ptr_r [2] ? _09883_ : _09880_;
  assign _09885_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [8] : \MSYNC_1r1w.synth.nz.mem[632] [8];
  assign _09886_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [8] : \MSYNC_1r1w.synth.nz.mem[634] [8];
  assign _09887_ = \bapg_rd.w_ptr_r [1] ? _09886_ : _09885_;
  assign _09888_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [8] : \MSYNC_1r1w.synth.nz.mem[636] [8];
  assign _09889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [8] : \MSYNC_1r1w.synth.nz.mem[638] [8];
  assign _09890_ = \bapg_rd.w_ptr_r [1] ? _09889_ : _09888_;
  assign _09891_ = \bapg_rd.w_ptr_r [2] ? _09890_ : _09887_;
  assign _09892_ = \bapg_rd.w_ptr_r [3] ? _09891_ : _09884_;
  assign _09893_ = \bapg_rd.w_ptr_r [4] ? _09892_ : _09877_;
  assign _09894_ = \bapg_rd.w_ptr_r [5] ? _09893_ : _09862_;
  assign _09895_ = \bapg_rd.w_ptr_r [6] ? _09894_ : _09831_;
  assign _09896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [8] : \MSYNC_1r1w.synth.nz.mem[640] [8];
  assign _09897_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [8] : \MSYNC_1r1w.synth.nz.mem[642] [8];
  assign _09898_ = \bapg_rd.w_ptr_r [1] ? _09897_ : _09896_;
  assign _09899_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [8] : \MSYNC_1r1w.synth.nz.mem[644] [8];
  assign _09900_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [8] : \MSYNC_1r1w.synth.nz.mem[646] [8];
  assign _09901_ = \bapg_rd.w_ptr_r [1] ? _09900_ : _09899_;
  assign _09902_ = \bapg_rd.w_ptr_r [2] ? _09901_ : _09898_;
  assign _09903_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [8] : \MSYNC_1r1w.synth.nz.mem[648] [8];
  assign _09904_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [8] : \MSYNC_1r1w.synth.nz.mem[650] [8];
  assign _09905_ = \bapg_rd.w_ptr_r [1] ? _09904_ : _09903_;
  assign _09906_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [8] : \MSYNC_1r1w.synth.nz.mem[652] [8];
  assign _09907_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [8] : \MSYNC_1r1w.synth.nz.mem[654] [8];
  assign _09908_ = \bapg_rd.w_ptr_r [1] ? _09907_ : _09906_;
  assign _09909_ = \bapg_rd.w_ptr_r [2] ? _09908_ : _09905_;
  assign _09910_ = \bapg_rd.w_ptr_r [3] ? _09909_ : _09902_;
  assign _09911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [8] : \MSYNC_1r1w.synth.nz.mem[656] [8];
  assign _09912_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [8] : \MSYNC_1r1w.synth.nz.mem[658] [8];
  assign _09913_ = \bapg_rd.w_ptr_r [1] ? _09912_ : _09911_;
  assign _09914_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [8] : \MSYNC_1r1w.synth.nz.mem[660] [8];
  assign _09915_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [8] : \MSYNC_1r1w.synth.nz.mem[662] [8];
  assign _09916_ = \bapg_rd.w_ptr_r [1] ? _09915_ : _09914_;
  assign _09917_ = \bapg_rd.w_ptr_r [2] ? _09916_ : _09913_;
  assign _09918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [8] : \MSYNC_1r1w.synth.nz.mem[664] [8];
  assign _09919_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [8] : \MSYNC_1r1w.synth.nz.mem[666] [8];
  assign _09920_ = \bapg_rd.w_ptr_r [1] ? _09919_ : _09918_;
  assign _09921_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [8] : \MSYNC_1r1w.synth.nz.mem[668] [8];
  assign _09922_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [8] : \MSYNC_1r1w.synth.nz.mem[670] [8];
  assign _09923_ = \bapg_rd.w_ptr_r [1] ? _09922_ : _09921_;
  assign _09924_ = \bapg_rd.w_ptr_r [2] ? _09923_ : _09920_;
  assign _09925_ = \bapg_rd.w_ptr_r [3] ? _09924_ : _09917_;
  assign _09926_ = \bapg_rd.w_ptr_r [4] ? _09925_ : _09910_;
  assign _09927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [8] : \MSYNC_1r1w.synth.nz.mem[672] [8];
  assign _09928_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [8] : \MSYNC_1r1w.synth.nz.mem[674] [8];
  assign _09929_ = \bapg_rd.w_ptr_r [1] ? _09928_ : _09927_;
  assign _09930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [8] : \MSYNC_1r1w.synth.nz.mem[676] [8];
  assign _09931_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [8] : \MSYNC_1r1w.synth.nz.mem[678] [8];
  assign _09932_ = \bapg_rd.w_ptr_r [1] ? _09931_ : _09930_;
  assign _09933_ = \bapg_rd.w_ptr_r [2] ? _09932_ : _09929_;
  assign _09934_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [8] : \MSYNC_1r1w.synth.nz.mem[680] [8];
  assign _09935_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [8] : \MSYNC_1r1w.synth.nz.mem[682] [8];
  assign _09936_ = \bapg_rd.w_ptr_r [1] ? _09935_ : _09934_;
  assign _09937_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [8] : \MSYNC_1r1w.synth.nz.mem[684] [8];
  assign _09938_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [8] : \MSYNC_1r1w.synth.nz.mem[686] [8];
  assign _09939_ = \bapg_rd.w_ptr_r [1] ? _09938_ : _09937_;
  assign _09940_ = \bapg_rd.w_ptr_r [2] ? _09939_ : _09936_;
  assign _09941_ = \bapg_rd.w_ptr_r [3] ? _09940_ : _09933_;
  assign _09942_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [8] : \MSYNC_1r1w.synth.nz.mem[688] [8];
  assign _09943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [8] : \MSYNC_1r1w.synth.nz.mem[690] [8];
  assign _09944_ = \bapg_rd.w_ptr_r [1] ? _09943_ : _09942_;
  assign _09945_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [8] : \MSYNC_1r1w.synth.nz.mem[692] [8];
  assign _09946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [8] : \MSYNC_1r1w.synth.nz.mem[694] [8];
  assign _09947_ = \bapg_rd.w_ptr_r [1] ? _09946_ : _09945_;
  assign _09948_ = \bapg_rd.w_ptr_r [2] ? _09947_ : _09944_;
  assign _09949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [8] : \MSYNC_1r1w.synth.nz.mem[696] [8];
  assign _09950_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [8] : \MSYNC_1r1w.synth.nz.mem[698] [8];
  assign _09951_ = \bapg_rd.w_ptr_r [1] ? _09950_ : _09949_;
  assign _09952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [8] : \MSYNC_1r1w.synth.nz.mem[700] [8];
  assign _09953_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [8] : \MSYNC_1r1w.synth.nz.mem[702] [8];
  assign _09954_ = \bapg_rd.w_ptr_r [1] ? _09953_ : _09952_;
  assign _09955_ = \bapg_rd.w_ptr_r [2] ? _09954_ : _09951_;
  assign _09956_ = \bapg_rd.w_ptr_r [3] ? _09955_ : _09948_;
  assign _09957_ = \bapg_rd.w_ptr_r [4] ? _09956_ : _09941_;
  assign _09958_ = \bapg_rd.w_ptr_r [5] ? _09957_ : _09926_;
  assign _09959_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [8] : \MSYNC_1r1w.synth.nz.mem[704] [8];
  assign _09960_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [8] : \MSYNC_1r1w.synth.nz.mem[706] [8];
  assign _09961_ = \bapg_rd.w_ptr_r [1] ? _09960_ : _09959_;
  assign _09962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [8] : \MSYNC_1r1w.synth.nz.mem[708] [8];
  assign _09963_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [8] : \MSYNC_1r1w.synth.nz.mem[710] [8];
  assign _09964_ = \bapg_rd.w_ptr_r [1] ? _09963_ : _09962_;
  assign _09965_ = \bapg_rd.w_ptr_r [2] ? _09964_ : _09961_;
  assign _09966_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [8] : \MSYNC_1r1w.synth.nz.mem[712] [8];
  assign _09967_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [8] : \MSYNC_1r1w.synth.nz.mem[714] [8];
  assign _09968_ = \bapg_rd.w_ptr_r [1] ? _09967_ : _09966_;
  assign _09969_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [8] : \MSYNC_1r1w.synth.nz.mem[716] [8];
  assign _09970_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [8] : \MSYNC_1r1w.synth.nz.mem[718] [8];
  assign _09971_ = \bapg_rd.w_ptr_r [1] ? _09970_ : _09969_;
  assign _09972_ = \bapg_rd.w_ptr_r [2] ? _09971_ : _09968_;
  assign _09973_ = \bapg_rd.w_ptr_r [3] ? _09972_ : _09965_;
  assign _09974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [8] : \MSYNC_1r1w.synth.nz.mem[720] [8];
  assign _09975_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [8] : \MSYNC_1r1w.synth.nz.mem[722] [8];
  assign _09976_ = \bapg_rd.w_ptr_r [1] ? _09975_ : _09974_;
  assign _09977_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [8] : \MSYNC_1r1w.synth.nz.mem[724] [8];
  assign _09978_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [8] : \MSYNC_1r1w.synth.nz.mem[726] [8];
  assign _09979_ = \bapg_rd.w_ptr_r [1] ? _09978_ : _09977_;
  assign _09980_ = \bapg_rd.w_ptr_r [2] ? _09979_ : _09976_;
  assign _09981_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [8] : \MSYNC_1r1w.synth.nz.mem[728] [8];
  assign _09982_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [8] : \MSYNC_1r1w.synth.nz.mem[730] [8];
  assign _09983_ = \bapg_rd.w_ptr_r [1] ? _09982_ : _09981_;
  assign _09984_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [8] : \MSYNC_1r1w.synth.nz.mem[732] [8];
  assign _09985_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [8] : \MSYNC_1r1w.synth.nz.mem[734] [8];
  assign _09986_ = \bapg_rd.w_ptr_r [1] ? _09985_ : _09984_;
  assign _09987_ = \bapg_rd.w_ptr_r [2] ? _09986_ : _09983_;
  assign _09988_ = \bapg_rd.w_ptr_r [3] ? _09987_ : _09980_;
  assign _09989_ = \bapg_rd.w_ptr_r [4] ? _09988_ : _09973_;
  assign _09990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [8] : \MSYNC_1r1w.synth.nz.mem[736] [8];
  assign _09991_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [8] : \MSYNC_1r1w.synth.nz.mem[738] [8];
  assign _09992_ = \bapg_rd.w_ptr_r [1] ? _09991_ : _09990_;
  assign _09993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [8] : \MSYNC_1r1w.synth.nz.mem[740] [8];
  assign _09994_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [8] : \MSYNC_1r1w.synth.nz.mem[742] [8];
  assign _09995_ = \bapg_rd.w_ptr_r [1] ? _09994_ : _09993_;
  assign _09996_ = \bapg_rd.w_ptr_r [2] ? _09995_ : _09992_;
  assign _09997_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [8] : \MSYNC_1r1w.synth.nz.mem[744] [8];
  assign _09998_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [8] : \MSYNC_1r1w.synth.nz.mem[746] [8];
  assign _09999_ = \bapg_rd.w_ptr_r [1] ? _09998_ : _09997_;
  assign _10000_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [8] : \MSYNC_1r1w.synth.nz.mem[748] [8];
  assign _10001_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [8] : \MSYNC_1r1w.synth.nz.mem[750] [8];
  assign _10002_ = \bapg_rd.w_ptr_r [1] ? _10001_ : _10000_;
  assign _10003_ = \bapg_rd.w_ptr_r [2] ? _10002_ : _09999_;
  assign _10004_ = \bapg_rd.w_ptr_r [3] ? _10003_ : _09996_;
  assign _10005_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [8] : \MSYNC_1r1w.synth.nz.mem[752] [8];
  assign _10006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [8] : \MSYNC_1r1w.synth.nz.mem[754] [8];
  assign _10007_ = \bapg_rd.w_ptr_r [1] ? _10006_ : _10005_;
  assign _10008_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [8] : \MSYNC_1r1w.synth.nz.mem[756] [8];
  assign _10009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [8] : \MSYNC_1r1w.synth.nz.mem[758] [8];
  assign _10010_ = \bapg_rd.w_ptr_r [1] ? _10009_ : _10008_;
  assign _10011_ = \bapg_rd.w_ptr_r [2] ? _10010_ : _10007_;
  assign _10012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [8] : \MSYNC_1r1w.synth.nz.mem[760] [8];
  assign _10013_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [8] : \MSYNC_1r1w.synth.nz.mem[762] [8];
  assign _10014_ = \bapg_rd.w_ptr_r [1] ? _10013_ : _10012_;
  assign _10015_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [8] : \MSYNC_1r1w.synth.nz.mem[764] [8];
  assign _10016_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [8] : \MSYNC_1r1w.synth.nz.mem[766] [8];
  assign _10017_ = \bapg_rd.w_ptr_r [1] ? _10016_ : _10015_;
  assign _10018_ = \bapg_rd.w_ptr_r [2] ? _10017_ : _10014_;
  assign _10019_ = \bapg_rd.w_ptr_r [3] ? _10018_ : _10011_;
  assign _10020_ = \bapg_rd.w_ptr_r [4] ? _10019_ : _10004_;
  assign _10021_ = \bapg_rd.w_ptr_r [5] ? _10020_ : _09989_;
  assign _10022_ = \bapg_rd.w_ptr_r [6] ? _10021_ : _09958_;
  assign _10023_ = \bapg_rd.w_ptr_r [7] ? _10022_ : _09895_;
  assign _10024_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [8] : \MSYNC_1r1w.synth.nz.mem[768] [8];
  assign _10025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [8] : \MSYNC_1r1w.synth.nz.mem[770] [8];
  assign _10026_ = \bapg_rd.w_ptr_r [1] ? _10025_ : _10024_;
  assign _10027_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [8] : \MSYNC_1r1w.synth.nz.mem[772] [8];
  assign _10028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [8] : \MSYNC_1r1w.synth.nz.mem[774] [8];
  assign _10029_ = \bapg_rd.w_ptr_r [1] ? _10028_ : _10027_;
  assign _10030_ = \bapg_rd.w_ptr_r [2] ? _10029_ : _10026_;
  assign _10031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [8] : \MSYNC_1r1w.synth.nz.mem[776] [8];
  assign _10032_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [8] : \MSYNC_1r1w.synth.nz.mem[778] [8];
  assign _10033_ = \bapg_rd.w_ptr_r [1] ? _10032_ : _10031_;
  assign _10034_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [8] : \MSYNC_1r1w.synth.nz.mem[780] [8];
  assign _10035_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [8] : \MSYNC_1r1w.synth.nz.mem[782] [8];
  assign _10036_ = \bapg_rd.w_ptr_r [1] ? _10035_ : _10034_;
  assign _10037_ = \bapg_rd.w_ptr_r [2] ? _10036_ : _10033_;
  assign _10038_ = \bapg_rd.w_ptr_r [3] ? _10037_ : _10030_;
  assign _10039_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [8] : \MSYNC_1r1w.synth.nz.mem[784] [8];
  assign _10040_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [8] : \MSYNC_1r1w.synth.nz.mem[786] [8];
  assign _10041_ = \bapg_rd.w_ptr_r [1] ? _10040_ : _10039_;
  assign _10042_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [8] : \MSYNC_1r1w.synth.nz.mem[788] [8];
  assign _10043_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [8] : \MSYNC_1r1w.synth.nz.mem[790] [8];
  assign _10044_ = \bapg_rd.w_ptr_r [1] ? _10043_ : _10042_;
  assign _10045_ = \bapg_rd.w_ptr_r [2] ? _10044_ : _10041_;
  assign _10046_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [8] : \MSYNC_1r1w.synth.nz.mem[792] [8];
  assign _10047_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [8] : \MSYNC_1r1w.synth.nz.mem[794] [8];
  assign _10048_ = \bapg_rd.w_ptr_r [1] ? _10047_ : _10046_;
  assign _10049_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [8] : \MSYNC_1r1w.synth.nz.mem[796] [8];
  assign _10050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [8] : \MSYNC_1r1w.synth.nz.mem[798] [8];
  assign _10051_ = \bapg_rd.w_ptr_r [1] ? _10050_ : _10049_;
  assign _10052_ = \bapg_rd.w_ptr_r [2] ? _10051_ : _10048_;
  assign _10053_ = \bapg_rd.w_ptr_r [3] ? _10052_ : _10045_;
  assign _10054_ = \bapg_rd.w_ptr_r [4] ? _10053_ : _10038_;
  assign _10055_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [8] : \MSYNC_1r1w.synth.nz.mem[800] [8];
  assign _10056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [8] : \MSYNC_1r1w.synth.nz.mem[802] [8];
  assign _10057_ = \bapg_rd.w_ptr_r [1] ? _10056_ : _10055_;
  assign _10058_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [8] : \MSYNC_1r1w.synth.nz.mem[804] [8];
  assign _10059_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [8] : \MSYNC_1r1w.synth.nz.mem[806] [8];
  assign _10060_ = \bapg_rd.w_ptr_r [1] ? _10059_ : _10058_;
  assign _10061_ = \bapg_rd.w_ptr_r [2] ? _10060_ : _10057_;
  assign _10062_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [8] : \MSYNC_1r1w.synth.nz.mem[808] [8];
  assign _10063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [8] : \MSYNC_1r1w.synth.nz.mem[810] [8];
  assign _10064_ = \bapg_rd.w_ptr_r [1] ? _10063_ : _10062_;
  assign _10065_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [8] : \MSYNC_1r1w.synth.nz.mem[812] [8];
  assign _10066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [8] : \MSYNC_1r1w.synth.nz.mem[814] [8];
  assign _10067_ = \bapg_rd.w_ptr_r [1] ? _10066_ : _10065_;
  assign _10068_ = \bapg_rd.w_ptr_r [2] ? _10067_ : _10064_;
  assign _10069_ = \bapg_rd.w_ptr_r [3] ? _10068_ : _10061_;
  assign _10070_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [8] : \MSYNC_1r1w.synth.nz.mem[816] [8];
  assign _10071_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [8] : \MSYNC_1r1w.synth.nz.mem[818] [8];
  assign _10072_ = \bapg_rd.w_ptr_r [1] ? _10071_ : _10070_;
  assign _10073_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [8] : \MSYNC_1r1w.synth.nz.mem[820] [8];
  assign _10074_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [8] : \MSYNC_1r1w.synth.nz.mem[822] [8];
  assign _10075_ = \bapg_rd.w_ptr_r [1] ? _10074_ : _10073_;
  assign _10076_ = \bapg_rd.w_ptr_r [2] ? _10075_ : _10072_;
  assign _10077_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [8] : \MSYNC_1r1w.synth.nz.mem[824] [8];
  assign _10078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [8] : \MSYNC_1r1w.synth.nz.mem[826] [8];
  assign _10079_ = \bapg_rd.w_ptr_r [1] ? _10078_ : _10077_;
  assign _10080_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [8] : \MSYNC_1r1w.synth.nz.mem[828] [8];
  assign _10081_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [8] : \MSYNC_1r1w.synth.nz.mem[830] [8];
  assign _10082_ = \bapg_rd.w_ptr_r [1] ? _10081_ : _10080_;
  assign _10083_ = \bapg_rd.w_ptr_r [2] ? _10082_ : _10079_;
  assign _10084_ = \bapg_rd.w_ptr_r [3] ? _10083_ : _10076_;
  assign _10085_ = \bapg_rd.w_ptr_r [4] ? _10084_ : _10069_;
  assign _10086_ = \bapg_rd.w_ptr_r [5] ? _10085_ : _10054_;
  assign _10087_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [8] : \MSYNC_1r1w.synth.nz.mem[832] [8];
  assign _10088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [8] : \MSYNC_1r1w.synth.nz.mem[834] [8];
  assign _10089_ = \bapg_rd.w_ptr_r [1] ? _10088_ : _10087_;
  assign _10090_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [8] : \MSYNC_1r1w.synth.nz.mem[836] [8];
  assign _10091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [8] : \MSYNC_1r1w.synth.nz.mem[838] [8];
  assign _10092_ = \bapg_rd.w_ptr_r [1] ? _10091_ : _10090_;
  assign _10093_ = \bapg_rd.w_ptr_r [2] ? _10092_ : _10089_;
  assign _10094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [8] : \MSYNC_1r1w.synth.nz.mem[840] [8];
  assign _10095_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [8] : \MSYNC_1r1w.synth.nz.mem[842] [8];
  assign _10096_ = \bapg_rd.w_ptr_r [1] ? _10095_ : _10094_;
  assign _10097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [8] : \MSYNC_1r1w.synth.nz.mem[844] [8];
  assign _10098_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [8] : \MSYNC_1r1w.synth.nz.mem[846] [8];
  assign _10099_ = \bapg_rd.w_ptr_r [1] ? _10098_ : _10097_;
  assign _10100_ = \bapg_rd.w_ptr_r [2] ? _10099_ : _10096_;
  assign _10101_ = \bapg_rd.w_ptr_r [3] ? _10100_ : _10093_;
  assign _10102_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [8] : \MSYNC_1r1w.synth.nz.mem[848] [8];
  assign _10103_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [8] : \MSYNC_1r1w.synth.nz.mem[850] [8];
  assign _10104_ = \bapg_rd.w_ptr_r [1] ? _10103_ : _10102_;
  assign _10105_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [8] : \MSYNC_1r1w.synth.nz.mem[852] [8];
  assign _10106_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [8] : \MSYNC_1r1w.synth.nz.mem[854] [8];
  assign _10107_ = \bapg_rd.w_ptr_r [1] ? _10106_ : _10105_;
  assign _10108_ = \bapg_rd.w_ptr_r [2] ? _10107_ : _10104_;
  assign _10109_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [8] : \MSYNC_1r1w.synth.nz.mem[856] [8];
  assign _10110_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [8] : \MSYNC_1r1w.synth.nz.mem[858] [8];
  assign _10111_ = \bapg_rd.w_ptr_r [1] ? _10110_ : _10109_;
  assign _10112_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [8] : \MSYNC_1r1w.synth.nz.mem[860] [8];
  assign _10113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [8] : \MSYNC_1r1w.synth.nz.mem[862] [8];
  assign _10114_ = \bapg_rd.w_ptr_r [1] ? _10113_ : _10112_;
  assign _10115_ = \bapg_rd.w_ptr_r [2] ? _10114_ : _10111_;
  assign _10116_ = \bapg_rd.w_ptr_r [3] ? _10115_ : _10108_;
  assign _10117_ = \bapg_rd.w_ptr_r [4] ? _10116_ : _10101_;
  assign _10118_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [8] : \MSYNC_1r1w.synth.nz.mem[864] [8];
  assign _10119_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [8] : \MSYNC_1r1w.synth.nz.mem[866] [8];
  assign _10120_ = \bapg_rd.w_ptr_r [1] ? _10119_ : _10118_;
  assign _10121_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [8] : \MSYNC_1r1w.synth.nz.mem[868] [8];
  assign _10122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [8] : \MSYNC_1r1w.synth.nz.mem[870] [8];
  assign _10123_ = \bapg_rd.w_ptr_r [1] ? _10122_ : _10121_;
  assign _10124_ = \bapg_rd.w_ptr_r [2] ? _10123_ : _10120_;
  assign _10125_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [8] : \MSYNC_1r1w.synth.nz.mem[872] [8];
  assign _10126_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [8] : \MSYNC_1r1w.synth.nz.mem[874] [8];
  assign _10127_ = \bapg_rd.w_ptr_r [1] ? _10126_ : _10125_;
  assign _10128_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [8] : \MSYNC_1r1w.synth.nz.mem[876] [8];
  assign _10129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [8] : \MSYNC_1r1w.synth.nz.mem[878] [8];
  assign _10130_ = \bapg_rd.w_ptr_r [1] ? _10129_ : _10128_;
  assign _10131_ = \bapg_rd.w_ptr_r [2] ? _10130_ : _10127_;
  assign _10132_ = \bapg_rd.w_ptr_r [3] ? _10131_ : _10124_;
  assign _10133_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [8] : \MSYNC_1r1w.synth.nz.mem[880] [8];
  assign _10134_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [8] : \MSYNC_1r1w.synth.nz.mem[882] [8];
  assign _10135_ = \bapg_rd.w_ptr_r [1] ? _10134_ : _10133_;
  assign _10136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [8] : \MSYNC_1r1w.synth.nz.mem[884] [8];
  assign _10137_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [8] : \MSYNC_1r1w.synth.nz.mem[886] [8];
  assign _10138_ = \bapg_rd.w_ptr_r [1] ? _10137_ : _10136_;
  assign _10139_ = \bapg_rd.w_ptr_r [2] ? _10138_ : _10135_;
  assign _10140_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [8] : \MSYNC_1r1w.synth.nz.mem[888] [8];
  assign _10141_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [8] : \MSYNC_1r1w.synth.nz.mem[890] [8];
  assign _10142_ = \bapg_rd.w_ptr_r [1] ? _10141_ : _10140_;
  assign _10143_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [8] : \MSYNC_1r1w.synth.nz.mem[892] [8];
  assign _10144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [8] : \MSYNC_1r1w.synth.nz.mem[894] [8];
  assign _10145_ = \bapg_rd.w_ptr_r [1] ? _10144_ : _10143_;
  assign _10146_ = \bapg_rd.w_ptr_r [2] ? _10145_ : _10142_;
  assign _10147_ = \bapg_rd.w_ptr_r [3] ? _10146_ : _10139_;
  assign _10148_ = \bapg_rd.w_ptr_r [4] ? _10147_ : _10132_;
  assign _10149_ = \bapg_rd.w_ptr_r [5] ? _10148_ : _10117_;
  assign _10150_ = \bapg_rd.w_ptr_r [6] ? _10149_ : _10086_;
  assign _10151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [8] : \MSYNC_1r1w.synth.nz.mem[896] [8];
  assign _10152_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [8] : \MSYNC_1r1w.synth.nz.mem[898] [8];
  assign _10153_ = \bapg_rd.w_ptr_r [1] ? _10152_ : _10151_;
  assign _10154_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [8] : \MSYNC_1r1w.synth.nz.mem[900] [8];
  assign _10155_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [8] : \MSYNC_1r1w.synth.nz.mem[902] [8];
  assign _10156_ = \bapg_rd.w_ptr_r [1] ? _10155_ : _10154_;
  assign _10157_ = \bapg_rd.w_ptr_r [2] ? _10156_ : _10153_;
  assign _10158_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [8] : \MSYNC_1r1w.synth.nz.mem[904] [8];
  assign _10159_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [8] : \MSYNC_1r1w.synth.nz.mem[906] [8];
  assign _10160_ = \bapg_rd.w_ptr_r [1] ? _10159_ : _10158_;
  assign _10161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [8] : \MSYNC_1r1w.synth.nz.mem[908] [8];
  assign _10162_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [8] : \MSYNC_1r1w.synth.nz.mem[910] [8];
  assign _10163_ = \bapg_rd.w_ptr_r [1] ? _10162_ : _10161_;
  assign _10164_ = \bapg_rd.w_ptr_r [2] ? _10163_ : _10160_;
  assign _10165_ = \bapg_rd.w_ptr_r [3] ? _10164_ : _10157_;
  assign _10166_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [8] : \MSYNC_1r1w.synth.nz.mem[912] [8];
  assign _10167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [8] : \MSYNC_1r1w.synth.nz.mem[914] [8];
  assign _10168_ = \bapg_rd.w_ptr_r [1] ? _10167_ : _10166_;
  assign _10169_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [8] : \MSYNC_1r1w.synth.nz.mem[916] [8];
  assign _10170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [8] : \MSYNC_1r1w.synth.nz.mem[918] [8];
  assign _10171_ = \bapg_rd.w_ptr_r [1] ? _10170_ : _10169_;
  assign _10172_ = \bapg_rd.w_ptr_r [2] ? _10171_ : _10168_;
  assign _10173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [8] : \MSYNC_1r1w.synth.nz.mem[920] [8];
  assign _10174_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [8] : \MSYNC_1r1w.synth.nz.mem[922] [8];
  assign _10175_ = \bapg_rd.w_ptr_r [1] ? _10174_ : _10173_;
  assign _10176_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [8] : \MSYNC_1r1w.synth.nz.mem[924] [8];
  assign _10177_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [8] : \MSYNC_1r1w.synth.nz.mem[926] [8];
  assign _10178_ = \bapg_rd.w_ptr_r [1] ? _10177_ : _10176_;
  assign _10179_ = \bapg_rd.w_ptr_r [2] ? _10178_ : _10175_;
  assign _10180_ = \bapg_rd.w_ptr_r [3] ? _10179_ : _10172_;
  assign _10181_ = \bapg_rd.w_ptr_r [4] ? _10180_ : _10165_;
  assign _10182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [8] : \MSYNC_1r1w.synth.nz.mem[928] [8];
  assign _10183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [8] : \MSYNC_1r1w.synth.nz.mem[930] [8];
  assign _10184_ = \bapg_rd.w_ptr_r [1] ? _10183_ : _10182_;
  assign _10185_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [8] : \MSYNC_1r1w.synth.nz.mem[932] [8];
  assign _10186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [8] : \MSYNC_1r1w.synth.nz.mem[934] [8];
  assign _10187_ = \bapg_rd.w_ptr_r [1] ? _10186_ : _10185_;
  assign _10188_ = \bapg_rd.w_ptr_r [2] ? _10187_ : _10184_;
  assign _10189_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [8] : \MSYNC_1r1w.synth.nz.mem[936] [8];
  assign _10190_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [8] : \MSYNC_1r1w.synth.nz.mem[938] [8];
  assign _10191_ = \bapg_rd.w_ptr_r [1] ? _10190_ : _10189_;
  assign _10192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [8] : \MSYNC_1r1w.synth.nz.mem[940] [8];
  assign _10193_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [8] : \MSYNC_1r1w.synth.nz.mem[942] [8];
  assign _10194_ = \bapg_rd.w_ptr_r [1] ? _10193_ : _10192_;
  assign _10195_ = \bapg_rd.w_ptr_r [2] ? _10194_ : _10191_;
  assign _10196_ = \bapg_rd.w_ptr_r [3] ? _10195_ : _10188_;
  assign _10197_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [8] : \MSYNC_1r1w.synth.nz.mem[944] [8];
  assign _10198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [8] : \MSYNC_1r1w.synth.nz.mem[946] [8];
  assign _10199_ = \bapg_rd.w_ptr_r [1] ? _10198_ : _10197_;
  assign _10200_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [8] : \MSYNC_1r1w.synth.nz.mem[948] [8];
  assign _10201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [8] : \MSYNC_1r1w.synth.nz.mem[950] [8];
  assign _10202_ = \bapg_rd.w_ptr_r [1] ? _10201_ : _10200_;
  assign _10203_ = \bapg_rd.w_ptr_r [2] ? _10202_ : _10199_;
  assign _10204_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [8] : \MSYNC_1r1w.synth.nz.mem[952] [8];
  assign _10205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [8] : \MSYNC_1r1w.synth.nz.mem[954] [8];
  assign _10206_ = \bapg_rd.w_ptr_r [1] ? _10205_ : _10204_;
  assign _10207_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [8] : \MSYNC_1r1w.synth.nz.mem[956] [8];
  assign _10208_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [8] : \MSYNC_1r1w.synth.nz.mem[958] [8];
  assign _10209_ = \bapg_rd.w_ptr_r [1] ? _10208_ : _10207_;
  assign _10210_ = \bapg_rd.w_ptr_r [2] ? _10209_ : _10206_;
  assign _10211_ = \bapg_rd.w_ptr_r [3] ? _10210_ : _10203_;
  assign _10212_ = \bapg_rd.w_ptr_r [4] ? _10211_ : _10196_;
  assign _10213_ = \bapg_rd.w_ptr_r [5] ? _10212_ : _10181_;
  assign _10214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [8] : \MSYNC_1r1w.synth.nz.mem[960] [8];
  assign _10215_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [8] : \MSYNC_1r1w.synth.nz.mem[962] [8];
  assign _10216_ = \bapg_rd.w_ptr_r [1] ? _10215_ : _10214_;
  assign _10217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [8] : \MSYNC_1r1w.synth.nz.mem[964] [8];
  assign _10218_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [8] : \MSYNC_1r1w.synth.nz.mem[966] [8];
  assign _10219_ = \bapg_rd.w_ptr_r [1] ? _10218_ : _10217_;
  assign _10220_ = \bapg_rd.w_ptr_r [2] ? _10219_ : _10216_;
  assign _10221_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [8] : \MSYNC_1r1w.synth.nz.mem[968] [8];
  assign _10222_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [8] : \MSYNC_1r1w.synth.nz.mem[970] [8];
  assign _10223_ = \bapg_rd.w_ptr_r [1] ? _10222_ : _10221_;
  assign _10224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [8] : \MSYNC_1r1w.synth.nz.mem[972] [8];
  assign _10225_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [8] : \MSYNC_1r1w.synth.nz.mem[974] [8];
  assign _10226_ = \bapg_rd.w_ptr_r [1] ? _10225_ : _10224_;
  assign _10227_ = \bapg_rd.w_ptr_r [2] ? _10226_ : _10223_;
  assign _10228_ = \bapg_rd.w_ptr_r [3] ? _10227_ : _10220_;
  assign _10229_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [8] : \MSYNC_1r1w.synth.nz.mem[976] [8];
  assign _10230_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [8] : \MSYNC_1r1w.synth.nz.mem[978] [8];
  assign _10231_ = \bapg_rd.w_ptr_r [1] ? _10230_ : _10229_;
  assign _10232_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [8] : \MSYNC_1r1w.synth.nz.mem[980] [8];
  assign _10233_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [8] : \MSYNC_1r1w.synth.nz.mem[982] [8];
  assign _10234_ = \bapg_rd.w_ptr_r [1] ? _10233_ : _10232_;
  assign _10235_ = \bapg_rd.w_ptr_r [2] ? _10234_ : _10231_;
  assign _10236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [8] : \MSYNC_1r1w.synth.nz.mem[984] [8];
  assign _10237_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [8] : \MSYNC_1r1w.synth.nz.mem[986] [8];
  assign _10238_ = \bapg_rd.w_ptr_r [1] ? _10237_ : _10236_;
  assign _10239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [8] : \MSYNC_1r1w.synth.nz.mem[988] [8];
  assign _10240_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [8] : \MSYNC_1r1w.synth.nz.mem[990] [8];
  assign _10241_ = \bapg_rd.w_ptr_r [1] ? _10240_ : _10239_;
  assign _10242_ = \bapg_rd.w_ptr_r [2] ? _10241_ : _10238_;
  assign _10243_ = \bapg_rd.w_ptr_r [3] ? _10242_ : _10235_;
  assign _10244_ = \bapg_rd.w_ptr_r [4] ? _10243_ : _10228_;
  assign _10245_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [8] : \MSYNC_1r1w.synth.nz.mem[992] [8];
  assign _10246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [8] : \MSYNC_1r1w.synth.nz.mem[994] [8];
  assign _10247_ = \bapg_rd.w_ptr_r [1] ? _10246_ : _10245_;
  assign _10248_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [8] : \MSYNC_1r1w.synth.nz.mem[996] [8];
  assign _10249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [8] : \MSYNC_1r1w.synth.nz.mem[998] [8];
  assign _10250_ = \bapg_rd.w_ptr_r [1] ? _10249_ : _10248_;
  assign _10251_ = \bapg_rd.w_ptr_r [2] ? _10250_ : _10247_;
  assign _10252_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [8] : \MSYNC_1r1w.synth.nz.mem[1000] [8];
  assign _10253_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [8] : \MSYNC_1r1w.synth.nz.mem[1002] [8];
  assign _10254_ = \bapg_rd.w_ptr_r [1] ? _10253_ : _10252_;
  assign _10255_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [8] : \MSYNC_1r1w.synth.nz.mem[1004] [8];
  assign _10256_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [8] : \MSYNC_1r1w.synth.nz.mem[1006] [8];
  assign _10257_ = \bapg_rd.w_ptr_r [1] ? _10256_ : _10255_;
  assign _10258_ = \bapg_rd.w_ptr_r [2] ? _10257_ : _10254_;
  assign _10259_ = \bapg_rd.w_ptr_r [3] ? _10258_ : _10251_;
  assign _10260_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [8] : \MSYNC_1r1w.synth.nz.mem[1008] [8];
  assign _10261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [8] : \MSYNC_1r1w.synth.nz.mem[1010] [8];
  assign _10262_ = \bapg_rd.w_ptr_r [1] ? _10261_ : _10260_;
  assign _10263_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [8] : \MSYNC_1r1w.synth.nz.mem[1012] [8];
  assign _10264_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [8] : \MSYNC_1r1w.synth.nz.mem[1014] [8];
  assign _10265_ = \bapg_rd.w_ptr_r [1] ? _10264_ : _10263_;
  assign _10266_ = \bapg_rd.w_ptr_r [2] ? _10265_ : _10262_;
  assign _10267_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [8] : \MSYNC_1r1w.synth.nz.mem[1016] [8];
  assign _10268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [8] : \MSYNC_1r1w.synth.nz.mem[1018] [8];
  assign _10269_ = \bapg_rd.w_ptr_r [1] ? _10268_ : _10267_;
  assign _10270_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [8] : \MSYNC_1r1w.synth.nz.mem[1020] [8];
  assign _10271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [8] : \MSYNC_1r1w.synth.nz.mem[1022] [8];
  assign _10272_ = \bapg_rd.w_ptr_r [1] ? _10271_ : _10270_;
  assign _10273_ = \bapg_rd.w_ptr_r [2] ? _10272_ : _10269_;
  assign _10274_ = \bapg_rd.w_ptr_r [3] ? _10273_ : _10266_;
  assign _10275_ = \bapg_rd.w_ptr_r [4] ? _10274_ : _10259_;
  assign _10276_ = \bapg_rd.w_ptr_r [5] ? _10275_ : _10244_;
  assign _10277_ = \bapg_rd.w_ptr_r [6] ? _10276_ : _10213_;
  assign _10278_ = \bapg_rd.w_ptr_r [7] ? _10277_ : _10150_;
  assign _10279_ = \bapg_rd.w_ptr_r [8] ? _10278_ : _10023_;
  assign r_data_o[8] = \bapg_rd.w_ptr_r [9] ? _10279_ : _09768_;
  assign _10280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [9] : \MSYNC_1r1w.synth.nz.mem[0] [9];
  assign _10281_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [9] : \MSYNC_1r1w.synth.nz.mem[2] [9];
  assign _10282_ = \bapg_rd.w_ptr_r [1] ? _10281_ : _10280_;
  assign _10283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [9] : \MSYNC_1r1w.synth.nz.mem[4] [9];
  assign _10284_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [9] : \MSYNC_1r1w.synth.nz.mem[6] [9];
  assign _10285_ = \bapg_rd.w_ptr_r [1] ? _10284_ : _10283_;
  assign _10286_ = \bapg_rd.w_ptr_r [2] ? _10285_ : _10282_;
  assign _10287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [9] : \MSYNC_1r1w.synth.nz.mem[8] [9];
  assign _10288_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [9] : \MSYNC_1r1w.synth.nz.mem[10] [9];
  assign _10289_ = \bapg_rd.w_ptr_r [1] ? _10288_ : _10287_;
  assign _10290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [9] : \MSYNC_1r1w.synth.nz.mem[12] [9];
  assign _10291_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [9] : \MSYNC_1r1w.synth.nz.mem[14] [9];
  assign _10292_ = \bapg_rd.w_ptr_r [1] ? _10291_ : _10290_;
  assign _10293_ = \bapg_rd.w_ptr_r [2] ? _10292_ : _10289_;
  assign _10294_ = \bapg_rd.w_ptr_r [3] ? _10293_ : _10286_;
  assign _10295_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [9] : \MSYNC_1r1w.synth.nz.mem[16] [9];
  assign _10296_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [9] : \MSYNC_1r1w.synth.nz.mem[18] [9];
  assign _10297_ = \bapg_rd.w_ptr_r [1] ? _10296_ : _10295_;
  assign _10298_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [9] : \MSYNC_1r1w.synth.nz.mem[20] [9];
  assign _10299_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [9] : \MSYNC_1r1w.synth.nz.mem[22] [9];
  assign _10300_ = \bapg_rd.w_ptr_r [1] ? _10299_ : _10298_;
  assign _10301_ = \bapg_rd.w_ptr_r [2] ? _10300_ : _10297_;
  assign _10302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [9] : \MSYNC_1r1w.synth.nz.mem[24] [9];
  assign _10303_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [9] : \MSYNC_1r1w.synth.nz.mem[26] [9];
  assign _10304_ = \bapg_rd.w_ptr_r [1] ? _10303_ : _10302_;
  assign _10305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [9] : \MSYNC_1r1w.synth.nz.mem[28] [9];
  assign _10306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [9] : \MSYNC_1r1w.synth.nz.mem[30] [9];
  assign _10307_ = \bapg_rd.w_ptr_r [1] ? _10306_ : _10305_;
  assign _10308_ = \bapg_rd.w_ptr_r [2] ? _10307_ : _10304_;
  assign _10309_ = \bapg_rd.w_ptr_r [3] ? _10308_ : _10301_;
  assign _10310_ = \bapg_rd.w_ptr_r [4] ? _10309_ : _10294_;
  assign _10311_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [9] : \MSYNC_1r1w.synth.nz.mem[32] [9];
  assign _10312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [9] : \MSYNC_1r1w.synth.nz.mem[34] [9];
  assign _10313_ = \bapg_rd.w_ptr_r [1] ? _10312_ : _10311_;
  assign _10314_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [9] : \MSYNC_1r1w.synth.nz.mem[36] [9];
  assign _10315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [9] : \MSYNC_1r1w.synth.nz.mem[38] [9];
  assign _10316_ = \bapg_rd.w_ptr_r [1] ? _10315_ : _10314_;
  assign _10317_ = \bapg_rd.w_ptr_r [2] ? _10316_ : _10313_;
  assign _10318_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [9] : \MSYNC_1r1w.synth.nz.mem[40] [9];
  assign _10319_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [9] : \MSYNC_1r1w.synth.nz.mem[42] [9];
  assign _10320_ = \bapg_rd.w_ptr_r [1] ? _10319_ : _10318_;
  assign _10321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [9] : \MSYNC_1r1w.synth.nz.mem[44] [9];
  assign _10322_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [9] : \MSYNC_1r1w.synth.nz.mem[46] [9];
  assign _10323_ = \bapg_rd.w_ptr_r [1] ? _10322_ : _10321_;
  assign _10324_ = \bapg_rd.w_ptr_r [2] ? _10323_ : _10320_;
  assign _10325_ = \bapg_rd.w_ptr_r [3] ? _10324_ : _10317_;
  assign _10326_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [9] : \MSYNC_1r1w.synth.nz.mem[48] [9];
  assign _10327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [9] : \MSYNC_1r1w.synth.nz.mem[50] [9];
  assign _10328_ = \bapg_rd.w_ptr_r [1] ? _10327_ : _10326_;
  assign _10329_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [9] : \MSYNC_1r1w.synth.nz.mem[52] [9];
  assign _10330_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [9] : \MSYNC_1r1w.synth.nz.mem[54] [9];
  assign _10331_ = \bapg_rd.w_ptr_r [1] ? _10330_ : _10329_;
  assign _10332_ = \bapg_rd.w_ptr_r [2] ? _10331_ : _10328_;
  assign _10333_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [9] : \MSYNC_1r1w.synth.nz.mem[56] [9];
  assign _10334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [9] : \MSYNC_1r1w.synth.nz.mem[58] [9];
  assign _10335_ = \bapg_rd.w_ptr_r [1] ? _10334_ : _10333_;
  assign _10336_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [9] : \MSYNC_1r1w.synth.nz.mem[60] [9];
  assign _10337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [9] : \MSYNC_1r1w.synth.nz.mem[62] [9];
  assign _10338_ = \bapg_rd.w_ptr_r [1] ? _10337_ : _10336_;
  assign _10339_ = \bapg_rd.w_ptr_r [2] ? _10338_ : _10335_;
  assign _10340_ = \bapg_rd.w_ptr_r [3] ? _10339_ : _10332_;
  assign _10341_ = \bapg_rd.w_ptr_r [4] ? _10340_ : _10325_;
  assign _10342_ = \bapg_rd.w_ptr_r [5] ? _10341_ : _10310_;
  assign _10343_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [9] : \MSYNC_1r1w.synth.nz.mem[64] [9];
  assign _10344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [9] : \MSYNC_1r1w.synth.nz.mem[66] [9];
  assign _10345_ = \bapg_rd.w_ptr_r [1] ? _10344_ : _10343_;
  assign _10346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [9] : \MSYNC_1r1w.synth.nz.mem[68] [9];
  assign _10347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [9] : \MSYNC_1r1w.synth.nz.mem[70] [9];
  assign _10348_ = \bapg_rd.w_ptr_r [1] ? _10347_ : _10346_;
  assign _10349_ = \bapg_rd.w_ptr_r [2] ? _10348_ : _10345_;
  assign _10350_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [9] : \MSYNC_1r1w.synth.nz.mem[72] [9];
  assign _10351_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [9] : \MSYNC_1r1w.synth.nz.mem[74] [9];
  assign _10352_ = \bapg_rd.w_ptr_r [1] ? _10351_ : _10350_;
  assign _10353_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [9] : \MSYNC_1r1w.synth.nz.mem[76] [9];
  assign _10354_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [9] : \MSYNC_1r1w.synth.nz.mem[78] [9];
  assign _10355_ = \bapg_rd.w_ptr_r [1] ? _10354_ : _10353_;
  assign _10356_ = \bapg_rd.w_ptr_r [2] ? _10355_ : _10352_;
  assign _10357_ = \bapg_rd.w_ptr_r [3] ? _10356_ : _10349_;
  assign _10358_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [9] : \MSYNC_1r1w.synth.nz.mem[80] [9];
  assign _10359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [9] : \MSYNC_1r1w.synth.nz.mem[82] [9];
  assign _10360_ = \bapg_rd.w_ptr_r [1] ? _10359_ : _10358_;
  assign _10361_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [9] : \MSYNC_1r1w.synth.nz.mem[84] [9];
  assign _10362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [9] : \MSYNC_1r1w.synth.nz.mem[86] [9];
  assign _10363_ = \bapg_rd.w_ptr_r [1] ? _10362_ : _10361_;
  assign _10364_ = \bapg_rd.w_ptr_r [2] ? _10363_ : _10360_;
  assign _10365_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [9] : \MSYNC_1r1w.synth.nz.mem[88] [9];
  assign _10366_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [9] : \MSYNC_1r1w.synth.nz.mem[90] [9];
  assign _10367_ = \bapg_rd.w_ptr_r [1] ? _10366_ : _10365_;
  assign _10368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [9] : \MSYNC_1r1w.synth.nz.mem[92] [9];
  assign _10369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [9] : \MSYNC_1r1w.synth.nz.mem[94] [9];
  assign _10370_ = \bapg_rd.w_ptr_r [1] ? _10369_ : _10368_;
  assign _10371_ = \bapg_rd.w_ptr_r [2] ? _10370_ : _10367_;
  assign _10372_ = \bapg_rd.w_ptr_r [3] ? _10371_ : _10364_;
  assign _10373_ = \bapg_rd.w_ptr_r [4] ? _10372_ : _10357_;
  assign _10374_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [9] : \MSYNC_1r1w.synth.nz.mem[96] [9];
  assign _10375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [9] : \MSYNC_1r1w.synth.nz.mem[98] [9];
  assign _10376_ = \bapg_rd.w_ptr_r [1] ? _10375_ : _10374_;
  assign _10377_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [9] : \MSYNC_1r1w.synth.nz.mem[100] [9];
  assign _10378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [9] : \MSYNC_1r1w.synth.nz.mem[102] [9];
  assign _10379_ = \bapg_rd.w_ptr_r [1] ? _10378_ : _10377_;
  assign _10380_ = \bapg_rd.w_ptr_r [2] ? _10379_ : _10376_;
  assign _10381_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [9] : \MSYNC_1r1w.synth.nz.mem[104] [9];
  assign _10382_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [9] : \MSYNC_1r1w.synth.nz.mem[106] [9];
  assign _10383_ = \bapg_rd.w_ptr_r [1] ? _10382_ : _10381_;
  assign _10384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [9] : \MSYNC_1r1w.synth.nz.mem[108] [9];
  assign _10385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [9] : \MSYNC_1r1w.synth.nz.mem[110] [9];
  assign _10386_ = \bapg_rd.w_ptr_r [1] ? _10385_ : _10384_;
  assign _10387_ = \bapg_rd.w_ptr_r [2] ? _10386_ : _10383_;
  assign _10388_ = \bapg_rd.w_ptr_r [3] ? _10387_ : _10380_;
  assign _10389_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [9] : \MSYNC_1r1w.synth.nz.mem[112] [9];
  assign _10390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [9] : \MSYNC_1r1w.synth.nz.mem[114] [9];
  assign _10391_ = \bapg_rd.w_ptr_r [1] ? _10390_ : _10389_;
  assign _10392_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [9] : \MSYNC_1r1w.synth.nz.mem[116] [9];
  assign _10393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [9] : \MSYNC_1r1w.synth.nz.mem[118] [9];
  assign _10394_ = \bapg_rd.w_ptr_r [1] ? _10393_ : _10392_;
  assign _10395_ = \bapg_rd.w_ptr_r [2] ? _10394_ : _10391_;
  assign _10396_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [9] : \MSYNC_1r1w.synth.nz.mem[120] [9];
  assign _10397_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [9] : \MSYNC_1r1w.synth.nz.mem[122] [9];
  assign _10398_ = \bapg_rd.w_ptr_r [1] ? _10397_ : _10396_;
  assign _10399_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [9] : \MSYNC_1r1w.synth.nz.mem[124] [9];
  assign _10400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [9] : \MSYNC_1r1w.synth.nz.mem[126] [9];
  assign _10401_ = \bapg_rd.w_ptr_r [1] ? _10400_ : _10399_;
  assign _10402_ = \bapg_rd.w_ptr_r [2] ? _10401_ : _10398_;
  assign _10403_ = \bapg_rd.w_ptr_r [3] ? _10402_ : _10395_;
  assign _10404_ = \bapg_rd.w_ptr_r [4] ? _10403_ : _10388_;
  assign _10405_ = \bapg_rd.w_ptr_r [5] ? _10404_ : _10373_;
  assign _10406_ = \bapg_rd.w_ptr_r [6] ? _10405_ : _10342_;
  assign _10407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [9] : \MSYNC_1r1w.synth.nz.mem[128] [9];
  assign _10408_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [9] : \MSYNC_1r1w.synth.nz.mem[130] [9];
  assign _10409_ = \bapg_rd.w_ptr_r [1] ? _10408_ : _10407_;
  assign _10410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [9] : \MSYNC_1r1w.synth.nz.mem[132] [9];
  assign _10411_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [9] : \MSYNC_1r1w.synth.nz.mem[134] [9];
  assign _10412_ = \bapg_rd.w_ptr_r [1] ? _10411_ : _10410_;
  assign _10413_ = \bapg_rd.w_ptr_r [2] ? _10412_ : _10409_;
  assign _10414_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [9] : \MSYNC_1r1w.synth.nz.mem[136] [9];
  assign _10415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [9] : \MSYNC_1r1w.synth.nz.mem[138] [9];
  assign _10416_ = \bapg_rd.w_ptr_r [1] ? _10415_ : _10414_;
  assign _10417_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [9] : \MSYNC_1r1w.synth.nz.mem[140] [9];
  assign _10418_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [9] : \MSYNC_1r1w.synth.nz.mem[142] [9];
  assign _10419_ = \bapg_rd.w_ptr_r [1] ? _10418_ : _10417_;
  assign _10420_ = \bapg_rd.w_ptr_r [2] ? _10419_ : _10416_;
  assign _10421_ = \bapg_rd.w_ptr_r [3] ? _10420_ : _10413_;
  assign _10422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [9] : \MSYNC_1r1w.synth.nz.mem[144] [9];
  assign _10423_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [9] : \MSYNC_1r1w.synth.nz.mem[146] [9];
  assign _10424_ = \bapg_rd.w_ptr_r [1] ? _10423_ : _10422_;
  assign _10425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [9] : \MSYNC_1r1w.synth.nz.mem[148] [9];
  assign _10426_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [9] : \MSYNC_1r1w.synth.nz.mem[150] [9];
  assign _10427_ = \bapg_rd.w_ptr_r [1] ? _10426_ : _10425_;
  assign _10428_ = \bapg_rd.w_ptr_r [2] ? _10427_ : _10424_;
  assign _10429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [9] : \MSYNC_1r1w.synth.nz.mem[152] [9];
  assign _10430_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [9] : \MSYNC_1r1w.synth.nz.mem[154] [9];
  assign _10431_ = \bapg_rd.w_ptr_r [1] ? _10430_ : _10429_;
  assign _10432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [9] : \MSYNC_1r1w.synth.nz.mem[156] [9];
  assign _10433_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [9] : \MSYNC_1r1w.synth.nz.mem[158] [9];
  assign _10434_ = \bapg_rd.w_ptr_r [1] ? _10433_ : _10432_;
  assign _10435_ = \bapg_rd.w_ptr_r [2] ? _10434_ : _10431_;
  assign _10436_ = \bapg_rd.w_ptr_r [3] ? _10435_ : _10428_;
  assign _10437_ = \bapg_rd.w_ptr_r [4] ? _10436_ : _10421_;
  assign _10438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [9] : \MSYNC_1r1w.synth.nz.mem[160] [9];
  assign _10439_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [9] : \MSYNC_1r1w.synth.nz.mem[162] [9];
  assign _10440_ = \bapg_rd.w_ptr_r [1] ? _10439_ : _10438_;
  assign _10441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [9] : \MSYNC_1r1w.synth.nz.mem[164] [9];
  assign _10442_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [9] : \MSYNC_1r1w.synth.nz.mem[166] [9];
  assign _10443_ = \bapg_rd.w_ptr_r [1] ? _10442_ : _10441_;
  assign _10444_ = \bapg_rd.w_ptr_r [2] ? _10443_ : _10440_;
  assign _10445_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [9] : \MSYNC_1r1w.synth.nz.mem[168] [9];
  assign _10446_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [9] : \MSYNC_1r1w.synth.nz.mem[170] [9];
  assign _10447_ = \bapg_rd.w_ptr_r [1] ? _10446_ : _10445_;
  assign _10448_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [9] : \MSYNC_1r1w.synth.nz.mem[172] [9];
  assign _10449_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [9] : \MSYNC_1r1w.synth.nz.mem[174] [9];
  assign _10450_ = \bapg_rd.w_ptr_r [1] ? _10449_ : _10448_;
  assign _10451_ = \bapg_rd.w_ptr_r [2] ? _10450_ : _10447_;
  assign _10452_ = \bapg_rd.w_ptr_r [3] ? _10451_ : _10444_;
  assign _10453_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [9] : \MSYNC_1r1w.synth.nz.mem[176] [9];
  assign _10454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [9] : \MSYNC_1r1w.synth.nz.mem[178] [9];
  assign _10455_ = \bapg_rd.w_ptr_r [1] ? _10454_ : _10453_;
  assign _10456_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [9] : \MSYNC_1r1w.synth.nz.mem[180] [9];
  assign _10457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [9] : \MSYNC_1r1w.synth.nz.mem[182] [9];
  assign _10458_ = \bapg_rd.w_ptr_r [1] ? _10457_ : _10456_;
  assign _10459_ = \bapg_rd.w_ptr_r [2] ? _10458_ : _10455_;
  assign _10460_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [9] : \MSYNC_1r1w.synth.nz.mem[184] [9];
  assign _10461_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [9] : \MSYNC_1r1w.synth.nz.mem[186] [9];
  assign _10462_ = \bapg_rd.w_ptr_r [1] ? _10461_ : _10460_;
  assign _10463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [9] : \MSYNC_1r1w.synth.nz.mem[188] [9];
  assign _10464_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [9] : \MSYNC_1r1w.synth.nz.mem[190] [9];
  assign _10465_ = \bapg_rd.w_ptr_r [1] ? _10464_ : _10463_;
  assign _10466_ = \bapg_rd.w_ptr_r [2] ? _10465_ : _10462_;
  assign _10467_ = \bapg_rd.w_ptr_r [3] ? _10466_ : _10459_;
  assign _10468_ = \bapg_rd.w_ptr_r [4] ? _10467_ : _10452_;
  assign _10469_ = \bapg_rd.w_ptr_r [5] ? _10468_ : _10437_;
  assign _10470_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [9] : \MSYNC_1r1w.synth.nz.mem[192] [9];
  assign _10471_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [9] : \MSYNC_1r1w.synth.nz.mem[194] [9];
  assign _10472_ = \bapg_rd.w_ptr_r [1] ? _10471_ : _10470_;
  assign _10473_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [9] : \MSYNC_1r1w.synth.nz.mem[196] [9];
  assign _10474_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [9] : \MSYNC_1r1w.synth.nz.mem[198] [9];
  assign _10475_ = \bapg_rd.w_ptr_r [1] ? _10474_ : _10473_;
  assign _10476_ = \bapg_rd.w_ptr_r [2] ? _10475_ : _10472_;
  assign _10477_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [9] : \MSYNC_1r1w.synth.nz.mem[200] [9];
  assign _10478_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [9] : \MSYNC_1r1w.synth.nz.mem[202] [9];
  assign _10479_ = \bapg_rd.w_ptr_r [1] ? _10478_ : _10477_;
  assign _10480_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [9] : \MSYNC_1r1w.synth.nz.mem[204] [9];
  assign _10481_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [9] : \MSYNC_1r1w.synth.nz.mem[206] [9];
  assign _10482_ = \bapg_rd.w_ptr_r [1] ? _10481_ : _10480_;
  assign _10483_ = \bapg_rd.w_ptr_r [2] ? _10482_ : _10479_;
  assign _10484_ = \bapg_rd.w_ptr_r [3] ? _10483_ : _10476_;
  assign _10485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [9] : \MSYNC_1r1w.synth.nz.mem[208] [9];
  assign _10486_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [9] : \MSYNC_1r1w.synth.nz.mem[210] [9];
  assign _10487_ = \bapg_rd.w_ptr_r [1] ? _10486_ : _10485_;
  assign _10488_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [9] : \MSYNC_1r1w.synth.nz.mem[212] [9];
  assign _10489_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [9] : \MSYNC_1r1w.synth.nz.mem[214] [9];
  assign _10490_ = \bapg_rd.w_ptr_r [1] ? _10489_ : _10488_;
  assign _10491_ = \bapg_rd.w_ptr_r [2] ? _10490_ : _10487_;
  assign _10492_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [9] : \MSYNC_1r1w.synth.nz.mem[216] [9];
  assign _10493_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [9] : \MSYNC_1r1w.synth.nz.mem[218] [9];
  assign _10494_ = \bapg_rd.w_ptr_r [1] ? _10493_ : _10492_;
  assign _10495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [9] : \MSYNC_1r1w.synth.nz.mem[220] [9];
  assign _10496_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [9] : \MSYNC_1r1w.synth.nz.mem[222] [9];
  assign _10497_ = \bapg_rd.w_ptr_r [1] ? _10496_ : _10495_;
  assign _10498_ = \bapg_rd.w_ptr_r [2] ? _10497_ : _10494_;
  assign _10499_ = \bapg_rd.w_ptr_r [3] ? _10498_ : _10491_;
  assign _10500_ = \bapg_rd.w_ptr_r [4] ? _10499_ : _10484_;
  assign _10501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [9] : \MSYNC_1r1w.synth.nz.mem[224] [9];
  assign _10502_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [9] : \MSYNC_1r1w.synth.nz.mem[226] [9];
  assign _10503_ = \bapg_rd.w_ptr_r [1] ? _10502_ : _10501_;
  assign _10504_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [9] : \MSYNC_1r1w.synth.nz.mem[228] [9];
  assign _10505_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [9] : \MSYNC_1r1w.synth.nz.mem[230] [9];
  assign _10506_ = \bapg_rd.w_ptr_r [1] ? _10505_ : _10504_;
  assign _10507_ = \bapg_rd.w_ptr_r [2] ? _10506_ : _10503_;
  assign _10508_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [9] : \MSYNC_1r1w.synth.nz.mem[232] [9];
  assign _10509_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [9] : \MSYNC_1r1w.synth.nz.mem[234] [9];
  assign _10510_ = \bapg_rd.w_ptr_r [1] ? _10509_ : _10508_;
  assign _10511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [9] : \MSYNC_1r1w.synth.nz.mem[236] [9];
  assign _10512_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [9] : \MSYNC_1r1w.synth.nz.mem[238] [9];
  assign _10513_ = \bapg_rd.w_ptr_r [1] ? _10512_ : _10511_;
  assign _10514_ = \bapg_rd.w_ptr_r [2] ? _10513_ : _10510_;
  assign _10515_ = \bapg_rd.w_ptr_r [3] ? _10514_ : _10507_;
  assign _10516_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [9] : \MSYNC_1r1w.synth.nz.mem[240] [9];
  assign _10517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [9] : \MSYNC_1r1w.synth.nz.mem[242] [9];
  assign _10518_ = \bapg_rd.w_ptr_r [1] ? _10517_ : _10516_;
  assign _10519_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [9] : \MSYNC_1r1w.synth.nz.mem[244] [9];
  assign _10520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [9] : \MSYNC_1r1w.synth.nz.mem[246] [9];
  assign _10521_ = \bapg_rd.w_ptr_r [1] ? _10520_ : _10519_;
  assign _10522_ = \bapg_rd.w_ptr_r [2] ? _10521_ : _10518_;
  assign _10523_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [9] : \MSYNC_1r1w.synth.nz.mem[248] [9];
  assign _10524_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [9] : \MSYNC_1r1w.synth.nz.mem[250] [9];
  assign _10525_ = \bapg_rd.w_ptr_r [1] ? _10524_ : _10523_;
  assign _10526_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [9] : \MSYNC_1r1w.synth.nz.mem[252] [9];
  assign _10527_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [9] : \MSYNC_1r1w.synth.nz.mem[254] [9];
  assign _10528_ = \bapg_rd.w_ptr_r [1] ? _10527_ : _10526_;
  assign _10529_ = \bapg_rd.w_ptr_r [2] ? _10528_ : _10525_;
  assign _10530_ = \bapg_rd.w_ptr_r [3] ? _10529_ : _10522_;
  assign _10531_ = \bapg_rd.w_ptr_r [4] ? _10530_ : _10515_;
  assign _10532_ = \bapg_rd.w_ptr_r [5] ? _10531_ : _10500_;
  assign _10533_ = \bapg_rd.w_ptr_r [6] ? _10532_ : _10469_;
  assign _10534_ = \bapg_rd.w_ptr_r [7] ? _10533_ : _10406_;
  assign _10535_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [9] : \MSYNC_1r1w.synth.nz.mem[256] [9];
  assign _10536_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [9] : \MSYNC_1r1w.synth.nz.mem[258] [9];
  assign _10537_ = \bapg_rd.w_ptr_r [1] ? _10536_ : _10535_;
  assign _10538_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [9] : \MSYNC_1r1w.synth.nz.mem[260] [9];
  assign _10539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [9] : \MSYNC_1r1w.synth.nz.mem[262] [9];
  assign _10540_ = \bapg_rd.w_ptr_r [1] ? _10539_ : _10538_;
  assign _10541_ = \bapg_rd.w_ptr_r [2] ? _10540_ : _10537_;
  assign _10542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [9] : \MSYNC_1r1w.synth.nz.mem[264] [9];
  assign _10543_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [9] : \MSYNC_1r1w.synth.nz.mem[266] [9];
  assign _10544_ = \bapg_rd.w_ptr_r [1] ? _10543_ : _10542_;
  assign _10545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [9] : \MSYNC_1r1w.synth.nz.mem[268] [9];
  assign _10546_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [9] : \MSYNC_1r1w.synth.nz.mem[270] [9];
  assign _10547_ = \bapg_rd.w_ptr_r [1] ? _10546_ : _10545_;
  assign _10548_ = \bapg_rd.w_ptr_r [2] ? _10547_ : _10544_;
  assign _10549_ = \bapg_rd.w_ptr_r [3] ? _10548_ : _10541_;
  assign _10550_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [9] : \MSYNC_1r1w.synth.nz.mem[272] [9];
  assign _10551_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [9] : \MSYNC_1r1w.synth.nz.mem[274] [9];
  assign _10552_ = \bapg_rd.w_ptr_r [1] ? _10551_ : _10550_;
  assign _10553_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [9] : \MSYNC_1r1w.synth.nz.mem[276] [9];
  assign _10554_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [9] : \MSYNC_1r1w.synth.nz.mem[278] [9];
  assign _10555_ = \bapg_rd.w_ptr_r [1] ? _10554_ : _10553_;
  assign _10556_ = \bapg_rd.w_ptr_r [2] ? _10555_ : _10552_;
  assign _10557_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [9] : \MSYNC_1r1w.synth.nz.mem[280] [9];
  assign _10558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [9] : \MSYNC_1r1w.synth.nz.mem[282] [9];
  assign _10559_ = \bapg_rd.w_ptr_r [1] ? _10558_ : _10557_;
  assign _10560_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [9] : \MSYNC_1r1w.synth.nz.mem[284] [9];
  assign _10561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [9] : \MSYNC_1r1w.synth.nz.mem[286] [9];
  assign _10562_ = \bapg_rd.w_ptr_r [1] ? _10561_ : _10560_;
  assign _10563_ = \bapg_rd.w_ptr_r [2] ? _10562_ : _10559_;
  assign _10564_ = \bapg_rd.w_ptr_r [3] ? _10563_ : _10556_;
  assign _10565_ = \bapg_rd.w_ptr_r [4] ? _10564_ : _10549_;
  assign _10566_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [9] : \MSYNC_1r1w.synth.nz.mem[288] [9];
  assign _10567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [9] : \MSYNC_1r1w.synth.nz.mem[290] [9];
  assign _10568_ = \bapg_rd.w_ptr_r [1] ? _10567_ : _10566_;
  assign _10569_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [9] : \MSYNC_1r1w.synth.nz.mem[292] [9];
  assign _10570_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [9] : \MSYNC_1r1w.synth.nz.mem[294] [9];
  assign _10571_ = \bapg_rd.w_ptr_r [1] ? _10570_ : _10569_;
  assign _10572_ = \bapg_rd.w_ptr_r [2] ? _10571_ : _10568_;
  assign _10573_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [9] : \MSYNC_1r1w.synth.nz.mem[296] [9];
  assign _10574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [9] : \MSYNC_1r1w.synth.nz.mem[298] [9];
  assign _10575_ = \bapg_rd.w_ptr_r [1] ? _10574_ : _10573_;
  assign _10576_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [9] : \MSYNC_1r1w.synth.nz.mem[300] [9];
  assign _10577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [9] : \MSYNC_1r1w.synth.nz.mem[302] [9];
  assign _10578_ = \bapg_rd.w_ptr_r [1] ? _10577_ : _10576_;
  assign _10579_ = \bapg_rd.w_ptr_r [2] ? _10578_ : _10575_;
  assign _10580_ = \bapg_rd.w_ptr_r [3] ? _10579_ : _10572_;
  assign _10581_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [9] : \MSYNC_1r1w.synth.nz.mem[304] [9];
  assign _10582_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [9] : \MSYNC_1r1w.synth.nz.mem[306] [9];
  assign _10583_ = \bapg_rd.w_ptr_r [1] ? _10582_ : _10581_;
  assign _10584_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [9] : \MSYNC_1r1w.synth.nz.mem[308] [9];
  assign _10585_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [9] : \MSYNC_1r1w.synth.nz.mem[310] [9];
  assign _10586_ = \bapg_rd.w_ptr_r [1] ? _10585_ : _10584_;
  assign _10587_ = \bapg_rd.w_ptr_r [2] ? _10586_ : _10583_;
  assign _10588_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [9] : \MSYNC_1r1w.synth.nz.mem[312] [9];
  assign _10589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [9] : \MSYNC_1r1w.synth.nz.mem[314] [9];
  assign _10590_ = \bapg_rd.w_ptr_r [1] ? _10589_ : _10588_;
  assign _10591_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [9] : \MSYNC_1r1w.synth.nz.mem[316] [9];
  assign _10592_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [9] : \MSYNC_1r1w.synth.nz.mem[318] [9];
  assign _10593_ = \bapg_rd.w_ptr_r [1] ? _10592_ : _10591_;
  assign _10594_ = \bapg_rd.w_ptr_r [2] ? _10593_ : _10590_;
  assign _10595_ = \bapg_rd.w_ptr_r [3] ? _10594_ : _10587_;
  assign _10596_ = \bapg_rd.w_ptr_r [4] ? _10595_ : _10580_;
  assign _10597_ = \bapg_rd.w_ptr_r [5] ? _10596_ : _10565_;
  assign _10598_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [9] : \MSYNC_1r1w.synth.nz.mem[320] [9];
  assign _10599_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [9] : \MSYNC_1r1w.synth.nz.mem[322] [9];
  assign _10600_ = \bapg_rd.w_ptr_r [1] ? _10599_ : _10598_;
  assign _10601_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [9] : \MSYNC_1r1w.synth.nz.mem[324] [9];
  assign _10602_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [9] : \MSYNC_1r1w.synth.nz.mem[326] [9];
  assign _10603_ = \bapg_rd.w_ptr_r [1] ? _10602_ : _10601_;
  assign _10604_ = \bapg_rd.w_ptr_r [2] ? _10603_ : _10600_;
  assign _10605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [9] : \MSYNC_1r1w.synth.nz.mem[328] [9];
  assign _10606_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [9] : \MSYNC_1r1w.synth.nz.mem[330] [9];
  assign _10607_ = \bapg_rd.w_ptr_r [1] ? _10606_ : _10605_;
  assign _10608_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [9] : \MSYNC_1r1w.synth.nz.mem[332] [9];
  assign _10609_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [9] : \MSYNC_1r1w.synth.nz.mem[334] [9];
  assign _10610_ = \bapg_rd.w_ptr_r [1] ? _10609_ : _10608_;
  assign _10611_ = \bapg_rd.w_ptr_r [2] ? _10610_ : _10607_;
  assign _10612_ = \bapg_rd.w_ptr_r [3] ? _10611_ : _10604_;
  assign _10613_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [9] : \MSYNC_1r1w.synth.nz.mem[336] [9];
  assign _10614_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [9] : \MSYNC_1r1w.synth.nz.mem[338] [9];
  assign _10615_ = \bapg_rd.w_ptr_r [1] ? _10614_ : _10613_;
  assign _10616_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [9] : \MSYNC_1r1w.synth.nz.mem[340] [9];
  assign _10617_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [9] : \MSYNC_1r1w.synth.nz.mem[342] [9];
  assign _10618_ = \bapg_rd.w_ptr_r [1] ? _10617_ : _10616_;
  assign _10619_ = \bapg_rd.w_ptr_r [2] ? _10618_ : _10615_;
  assign _10620_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [9] : \MSYNC_1r1w.synth.nz.mem[344] [9];
  assign _10621_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [9] : \MSYNC_1r1w.synth.nz.mem[346] [9];
  assign _10622_ = \bapg_rd.w_ptr_r [1] ? _10621_ : _10620_;
  assign _10623_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [9] : \MSYNC_1r1w.synth.nz.mem[348] [9];
  assign _10624_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [9] : \MSYNC_1r1w.synth.nz.mem[350] [9];
  assign _10625_ = \bapg_rd.w_ptr_r [1] ? _10624_ : _10623_;
  assign _10626_ = \bapg_rd.w_ptr_r [2] ? _10625_ : _10622_;
  assign _10627_ = \bapg_rd.w_ptr_r [3] ? _10626_ : _10619_;
  assign _10628_ = \bapg_rd.w_ptr_r [4] ? _10627_ : _10612_;
  assign _10629_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [9] : \MSYNC_1r1w.synth.nz.mem[352] [9];
  assign _10630_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [9] : \MSYNC_1r1w.synth.nz.mem[354] [9];
  assign _10631_ = \bapg_rd.w_ptr_r [1] ? _10630_ : _10629_;
  assign _10632_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [9] : \MSYNC_1r1w.synth.nz.mem[356] [9];
  assign _10633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [9] : \MSYNC_1r1w.synth.nz.mem[358] [9];
  assign _10634_ = \bapg_rd.w_ptr_r [1] ? _10633_ : _10632_;
  assign _10635_ = \bapg_rd.w_ptr_r [2] ? _10634_ : _10631_;
  assign _10636_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [9] : \MSYNC_1r1w.synth.nz.mem[360] [9];
  assign _10637_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [9] : \MSYNC_1r1w.synth.nz.mem[362] [9];
  assign _10638_ = \bapg_rd.w_ptr_r [1] ? _10637_ : _10636_;
  assign _10639_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [9] : \MSYNC_1r1w.synth.nz.mem[364] [9];
  assign _10640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [9] : \MSYNC_1r1w.synth.nz.mem[366] [9];
  assign _10641_ = \bapg_rd.w_ptr_r [1] ? _10640_ : _10639_;
  assign _10642_ = \bapg_rd.w_ptr_r [2] ? _10641_ : _10638_;
  assign _10643_ = \bapg_rd.w_ptr_r [3] ? _10642_ : _10635_;
  assign _10644_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [9] : \MSYNC_1r1w.synth.nz.mem[368] [9];
  assign _10645_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [9] : \MSYNC_1r1w.synth.nz.mem[370] [9];
  assign _10646_ = \bapg_rd.w_ptr_r [1] ? _10645_ : _10644_;
  assign _10647_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [9] : \MSYNC_1r1w.synth.nz.mem[372] [9];
  assign _10648_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [9] : \MSYNC_1r1w.synth.nz.mem[374] [9];
  assign _10649_ = \bapg_rd.w_ptr_r [1] ? _10648_ : _10647_;
  assign _10650_ = \bapg_rd.w_ptr_r [2] ? _10649_ : _10646_;
  assign _10651_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [9] : \MSYNC_1r1w.synth.nz.mem[376] [9];
  assign _10652_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [9] : \MSYNC_1r1w.synth.nz.mem[378] [9];
  assign _10653_ = \bapg_rd.w_ptr_r [1] ? _10652_ : _10651_;
  assign _10654_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [9] : \MSYNC_1r1w.synth.nz.mem[380] [9];
  assign _10655_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [9] : \MSYNC_1r1w.synth.nz.mem[382] [9];
  assign _10656_ = \bapg_rd.w_ptr_r [1] ? _10655_ : _10654_;
  assign _10657_ = \bapg_rd.w_ptr_r [2] ? _10656_ : _10653_;
  assign _10658_ = \bapg_rd.w_ptr_r [3] ? _10657_ : _10650_;
  assign _10659_ = \bapg_rd.w_ptr_r [4] ? _10658_ : _10643_;
  assign _10660_ = \bapg_rd.w_ptr_r [5] ? _10659_ : _10628_;
  assign _10661_ = \bapg_rd.w_ptr_r [6] ? _10660_ : _10597_;
  assign _10662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [9] : \MSYNC_1r1w.synth.nz.mem[384] [9];
  assign _10663_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [9] : \MSYNC_1r1w.synth.nz.mem[386] [9];
  assign _10664_ = \bapg_rd.w_ptr_r [1] ? _10663_ : _10662_;
  assign _10665_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [9] : \MSYNC_1r1w.synth.nz.mem[388] [9];
  assign _10666_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [9] : \MSYNC_1r1w.synth.nz.mem[390] [9];
  assign _10667_ = \bapg_rd.w_ptr_r [1] ? _10666_ : _10665_;
  assign _10668_ = \bapg_rd.w_ptr_r [2] ? _10667_ : _10664_;
  assign _10669_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [9] : \MSYNC_1r1w.synth.nz.mem[392] [9];
  assign _10670_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [9] : \MSYNC_1r1w.synth.nz.mem[394] [9];
  assign _10671_ = \bapg_rd.w_ptr_r [1] ? _10670_ : _10669_;
  assign _10672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [9] : \MSYNC_1r1w.synth.nz.mem[396] [9];
  assign _10673_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [9] : \MSYNC_1r1w.synth.nz.mem[398] [9];
  assign _10674_ = \bapg_rd.w_ptr_r [1] ? _10673_ : _10672_;
  assign _10675_ = \bapg_rd.w_ptr_r [2] ? _10674_ : _10671_;
  assign _10676_ = \bapg_rd.w_ptr_r [3] ? _10675_ : _10668_;
  assign _10677_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [9] : \MSYNC_1r1w.synth.nz.mem[400] [9];
  assign _10678_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [9] : \MSYNC_1r1w.synth.nz.mem[402] [9];
  assign _10679_ = \bapg_rd.w_ptr_r [1] ? _10678_ : _10677_;
  assign _10680_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [9] : \MSYNC_1r1w.synth.nz.mem[404] [9];
  assign _10681_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [9] : \MSYNC_1r1w.synth.nz.mem[406] [9];
  assign _10682_ = \bapg_rd.w_ptr_r [1] ? _10681_ : _10680_;
  assign _10683_ = \bapg_rd.w_ptr_r [2] ? _10682_ : _10679_;
  assign _10684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [9] : \MSYNC_1r1w.synth.nz.mem[408] [9];
  assign _10685_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [9] : \MSYNC_1r1w.synth.nz.mem[410] [9];
  assign _10686_ = \bapg_rd.w_ptr_r [1] ? _10685_ : _10684_;
  assign _10687_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [9] : \MSYNC_1r1w.synth.nz.mem[412] [9];
  assign _10688_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [9] : \MSYNC_1r1w.synth.nz.mem[414] [9];
  assign _10689_ = \bapg_rd.w_ptr_r [1] ? _10688_ : _10687_;
  assign _10690_ = \bapg_rd.w_ptr_r [2] ? _10689_ : _10686_;
  assign _10691_ = \bapg_rd.w_ptr_r [3] ? _10690_ : _10683_;
  assign _10692_ = \bapg_rd.w_ptr_r [4] ? _10691_ : _10676_;
  assign _10693_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [9] : \MSYNC_1r1w.synth.nz.mem[416] [9];
  assign _10694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [9] : \MSYNC_1r1w.synth.nz.mem[418] [9];
  assign _10695_ = \bapg_rd.w_ptr_r [1] ? _10694_ : _10693_;
  assign _10696_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [9] : \MSYNC_1r1w.synth.nz.mem[420] [9];
  assign _10697_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [9] : \MSYNC_1r1w.synth.nz.mem[422] [9];
  assign _10698_ = \bapg_rd.w_ptr_r [1] ? _10697_ : _10696_;
  assign _10699_ = \bapg_rd.w_ptr_r [2] ? _10698_ : _10695_;
  assign _10700_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [9] : \MSYNC_1r1w.synth.nz.mem[424] [9];
  assign _10701_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [9] : \MSYNC_1r1w.synth.nz.mem[426] [9];
  assign _10702_ = \bapg_rd.w_ptr_r [1] ? _10701_ : _10700_;
  assign _10703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [9] : \MSYNC_1r1w.synth.nz.mem[428] [9];
  assign _10704_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [9] : \MSYNC_1r1w.synth.nz.mem[430] [9];
  assign _10705_ = \bapg_rd.w_ptr_r [1] ? _10704_ : _10703_;
  assign _10706_ = \bapg_rd.w_ptr_r [2] ? _10705_ : _10702_;
  assign _10707_ = \bapg_rd.w_ptr_r [3] ? _10706_ : _10699_;
  assign _10708_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [9] : \MSYNC_1r1w.synth.nz.mem[432] [9];
  assign _10709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [9] : \MSYNC_1r1w.synth.nz.mem[434] [9];
  assign _10710_ = \bapg_rd.w_ptr_r [1] ? _10709_ : _10708_;
  assign _10711_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [9] : \MSYNC_1r1w.synth.nz.mem[436] [9];
  assign _10712_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [9] : \MSYNC_1r1w.synth.nz.mem[438] [9];
  assign _10713_ = \bapg_rd.w_ptr_r [1] ? _10712_ : _10711_;
  assign _10714_ = \bapg_rd.w_ptr_r [2] ? _10713_ : _10710_;
  assign _10715_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [9] : \MSYNC_1r1w.synth.nz.mem[440] [9];
  assign _10716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [9] : \MSYNC_1r1w.synth.nz.mem[442] [9];
  assign _10717_ = \bapg_rd.w_ptr_r [1] ? _10716_ : _10715_;
  assign _10718_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [9] : \MSYNC_1r1w.synth.nz.mem[444] [9];
  assign _10719_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [9] : \MSYNC_1r1w.synth.nz.mem[446] [9];
  assign _10720_ = \bapg_rd.w_ptr_r [1] ? _10719_ : _10718_;
  assign _10721_ = \bapg_rd.w_ptr_r [2] ? _10720_ : _10717_;
  assign _10722_ = \bapg_rd.w_ptr_r [3] ? _10721_ : _10714_;
  assign _10723_ = \bapg_rd.w_ptr_r [4] ? _10722_ : _10707_;
  assign _10724_ = \bapg_rd.w_ptr_r [5] ? _10723_ : _10692_;
  assign _10725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [9] : \MSYNC_1r1w.synth.nz.mem[448] [9];
  assign _10726_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [9] : \MSYNC_1r1w.synth.nz.mem[450] [9];
  assign _10727_ = \bapg_rd.w_ptr_r [1] ? _10726_ : _10725_;
  assign _10728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [9] : \MSYNC_1r1w.synth.nz.mem[452] [9];
  assign _10729_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [9] : \MSYNC_1r1w.synth.nz.mem[454] [9];
  assign _10730_ = \bapg_rd.w_ptr_r [1] ? _10729_ : _10728_;
  assign _10731_ = \bapg_rd.w_ptr_r [2] ? _10730_ : _10727_;
  assign _10732_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [9] : \MSYNC_1r1w.synth.nz.mem[456] [9];
  assign _10733_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [9] : \MSYNC_1r1w.synth.nz.mem[458] [9];
  assign _10734_ = \bapg_rd.w_ptr_r [1] ? _10733_ : _10732_;
  assign _10735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [9] : \MSYNC_1r1w.synth.nz.mem[460] [9];
  assign _10736_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [9] : \MSYNC_1r1w.synth.nz.mem[462] [9];
  assign _10737_ = \bapg_rd.w_ptr_r [1] ? _10736_ : _10735_;
  assign _10738_ = \bapg_rd.w_ptr_r [2] ? _10737_ : _10734_;
  assign _10739_ = \bapg_rd.w_ptr_r [3] ? _10738_ : _10731_;
  assign _10740_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [9] : \MSYNC_1r1w.synth.nz.mem[464] [9];
  assign _10741_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [9] : \MSYNC_1r1w.synth.nz.mem[466] [9];
  assign _10742_ = \bapg_rd.w_ptr_r [1] ? _10741_ : _10740_;
  assign _10743_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [9] : \MSYNC_1r1w.synth.nz.mem[468] [9];
  assign _10744_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [9] : \MSYNC_1r1w.synth.nz.mem[470] [9];
  assign _10745_ = \bapg_rd.w_ptr_r [1] ? _10744_ : _10743_;
  assign _10746_ = \bapg_rd.w_ptr_r [2] ? _10745_ : _10742_;
  assign _10747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [9] : \MSYNC_1r1w.synth.nz.mem[472] [9];
  assign _10748_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [9] : \MSYNC_1r1w.synth.nz.mem[474] [9];
  assign _10749_ = \bapg_rd.w_ptr_r [1] ? _10748_ : _10747_;
  assign _10750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [9] : \MSYNC_1r1w.synth.nz.mem[476] [9];
  assign _10751_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [9] : \MSYNC_1r1w.synth.nz.mem[478] [9];
  assign _10752_ = \bapg_rd.w_ptr_r [1] ? _10751_ : _10750_;
  assign _10753_ = \bapg_rd.w_ptr_r [2] ? _10752_ : _10749_;
  assign _10754_ = \bapg_rd.w_ptr_r [3] ? _10753_ : _10746_;
  assign _10755_ = \bapg_rd.w_ptr_r [4] ? _10754_ : _10739_;
  assign _10756_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [9] : \MSYNC_1r1w.synth.nz.mem[480] [9];
  assign _10757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [9] : \MSYNC_1r1w.synth.nz.mem[482] [9];
  assign _10758_ = \bapg_rd.w_ptr_r [1] ? _10757_ : _10756_;
  assign _10759_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [9] : \MSYNC_1r1w.synth.nz.mem[484] [9];
  assign _10760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [9] : \MSYNC_1r1w.synth.nz.mem[486] [9];
  assign _10761_ = \bapg_rd.w_ptr_r [1] ? _10760_ : _10759_;
  assign _10762_ = \bapg_rd.w_ptr_r [2] ? _10761_ : _10758_;
  assign _10763_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [9] : \MSYNC_1r1w.synth.nz.mem[488] [9];
  assign _10764_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [9] : \MSYNC_1r1w.synth.nz.mem[490] [9];
  assign _10765_ = \bapg_rd.w_ptr_r [1] ? _10764_ : _10763_;
  assign _10766_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [9] : \MSYNC_1r1w.synth.nz.mem[492] [9];
  assign _10767_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [9] : \MSYNC_1r1w.synth.nz.mem[494] [9];
  assign _10768_ = \bapg_rd.w_ptr_r [1] ? _10767_ : _10766_;
  assign _10769_ = \bapg_rd.w_ptr_r [2] ? _10768_ : _10765_;
  assign _10770_ = \bapg_rd.w_ptr_r [3] ? _10769_ : _10762_;
  assign _10771_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [9] : \MSYNC_1r1w.synth.nz.mem[496] [9];
  assign _10772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [9] : \MSYNC_1r1w.synth.nz.mem[498] [9];
  assign _10773_ = \bapg_rd.w_ptr_r [1] ? _10772_ : _10771_;
  assign _10774_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [9] : \MSYNC_1r1w.synth.nz.mem[500] [9];
  assign _10775_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [9] : \MSYNC_1r1w.synth.nz.mem[502] [9];
  assign _10776_ = \bapg_rd.w_ptr_r [1] ? _10775_ : _10774_;
  assign _10777_ = \bapg_rd.w_ptr_r [2] ? _10776_ : _10773_;
  assign _10778_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [9] : \MSYNC_1r1w.synth.nz.mem[504] [9];
  assign _10779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [9] : \MSYNC_1r1w.synth.nz.mem[506] [9];
  assign _10780_ = \bapg_rd.w_ptr_r [1] ? _10779_ : _10778_;
  assign _10781_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [9] : \MSYNC_1r1w.synth.nz.mem[508] [9];
  assign _10782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [9] : \MSYNC_1r1w.synth.nz.mem[510] [9];
  assign _10783_ = \bapg_rd.w_ptr_r [1] ? _10782_ : _10781_;
  assign _10784_ = \bapg_rd.w_ptr_r [2] ? _10783_ : _10780_;
  assign _10785_ = \bapg_rd.w_ptr_r [3] ? _10784_ : _10777_;
  assign _10786_ = \bapg_rd.w_ptr_r [4] ? _10785_ : _10770_;
  assign _10787_ = \bapg_rd.w_ptr_r [5] ? _10786_ : _10755_;
  assign _10788_ = \bapg_rd.w_ptr_r [6] ? _10787_ : _10724_;
  assign _10789_ = \bapg_rd.w_ptr_r [7] ? _10788_ : _10661_;
  assign _10790_ = \bapg_rd.w_ptr_r [8] ? _10789_ : _10534_;
  assign _10791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [9] : \MSYNC_1r1w.synth.nz.mem[512] [9];
  assign _10792_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [9] : \MSYNC_1r1w.synth.nz.mem[514] [9];
  assign _10793_ = \bapg_rd.w_ptr_r [1] ? _10792_ : _10791_;
  assign _10794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [9] : \MSYNC_1r1w.synth.nz.mem[516] [9];
  assign _10795_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [9] : \MSYNC_1r1w.synth.nz.mem[518] [9];
  assign _10796_ = \bapg_rd.w_ptr_r [1] ? _10795_ : _10794_;
  assign _10797_ = \bapg_rd.w_ptr_r [2] ? _10796_ : _10793_;
  assign _10798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [9] : \MSYNC_1r1w.synth.nz.mem[520] [9];
  assign _10799_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [9] : \MSYNC_1r1w.synth.nz.mem[522] [9];
  assign _10800_ = \bapg_rd.w_ptr_r [1] ? _10799_ : _10798_;
  assign _10801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [9] : \MSYNC_1r1w.synth.nz.mem[524] [9];
  assign _10802_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [9] : \MSYNC_1r1w.synth.nz.mem[526] [9];
  assign _10803_ = \bapg_rd.w_ptr_r [1] ? _10802_ : _10801_;
  assign _10804_ = \bapg_rd.w_ptr_r [2] ? _10803_ : _10800_;
  assign _10805_ = \bapg_rd.w_ptr_r [3] ? _10804_ : _10797_;
  assign _10806_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [9] : \MSYNC_1r1w.synth.nz.mem[528] [9];
  assign _10807_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [9] : \MSYNC_1r1w.synth.nz.mem[530] [9];
  assign _10808_ = \bapg_rd.w_ptr_r [1] ? _10807_ : _10806_;
  assign _10809_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [9] : \MSYNC_1r1w.synth.nz.mem[532] [9];
  assign _10810_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [9] : \MSYNC_1r1w.synth.nz.mem[534] [9];
  assign _10811_ = \bapg_rd.w_ptr_r [1] ? _10810_ : _10809_;
  assign _10812_ = \bapg_rd.w_ptr_r [2] ? _10811_ : _10808_;
  assign _10813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [9] : \MSYNC_1r1w.synth.nz.mem[536] [9];
  assign _10814_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [9] : \MSYNC_1r1w.synth.nz.mem[538] [9];
  assign _10815_ = \bapg_rd.w_ptr_r [1] ? _10814_ : _10813_;
  assign _10816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [9] : \MSYNC_1r1w.synth.nz.mem[540] [9];
  assign _10817_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [9] : \MSYNC_1r1w.synth.nz.mem[542] [9];
  assign _10818_ = \bapg_rd.w_ptr_r [1] ? _10817_ : _10816_;
  assign _10819_ = \bapg_rd.w_ptr_r [2] ? _10818_ : _10815_;
  assign _10820_ = \bapg_rd.w_ptr_r [3] ? _10819_ : _10812_;
  assign _10821_ = \bapg_rd.w_ptr_r [4] ? _10820_ : _10805_;
  assign _10822_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [9] : \MSYNC_1r1w.synth.nz.mem[544] [9];
  assign _10823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [9] : \MSYNC_1r1w.synth.nz.mem[546] [9];
  assign _10824_ = \bapg_rd.w_ptr_r [1] ? _10823_ : _10822_;
  assign _10825_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [9] : \MSYNC_1r1w.synth.nz.mem[548] [9];
  assign _10826_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [9] : \MSYNC_1r1w.synth.nz.mem[550] [9];
  assign _10827_ = \bapg_rd.w_ptr_r [1] ? _10826_ : _10825_;
  assign _10828_ = \bapg_rd.w_ptr_r [2] ? _10827_ : _10824_;
  assign _10829_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [9] : \MSYNC_1r1w.synth.nz.mem[552] [9];
  assign _10830_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [9] : \MSYNC_1r1w.synth.nz.mem[554] [9];
  assign _10831_ = \bapg_rd.w_ptr_r [1] ? _10830_ : _10829_;
  assign _10832_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [9] : \MSYNC_1r1w.synth.nz.mem[556] [9];
  assign _10833_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [9] : \MSYNC_1r1w.synth.nz.mem[558] [9];
  assign _10834_ = \bapg_rd.w_ptr_r [1] ? _10833_ : _10832_;
  assign _10835_ = \bapg_rd.w_ptr_r [2] ? _10834_ : _10831_;
  assign _10836_ = \bapg_rd.w_ptr_r [3] ? _10835_ : _10828_;
  assign _10837_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [9] : \MSYNC_1r1w.synth.nz.mem[560] [9];
  assign _10838_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [9] : \MSYNC_1r1w.synth.nz.mem[562] [9];
  assign _10839_ = \bapg_rd.w_ptr_r [1] ? _10838_ : _10837_;
  assign _10840_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [9] : \MSYNC_1r1w.synth.nz.mem[564] [9];
  assign _10841_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [9] : \MSYNC_1r1w.synth.nz.mem[566] [9];
  assign _10842_ = \bapg_rd.w_ptr_r [1] ? _10841_ : _10840_;
  assign _10843_ = \bapg_rd.w_ptr_r [2] ? _10842_ : _10839_;
  assign _10844_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [9] : \MSYNC_1r1w.synth.nz.mem[568] [9];
  assign _10845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [9] : \MSYNC_1r1w.synth.nz.mem[570] [9];
  assign _10846_ = \bapg_rd.w_ptr_r [1] ? _10845_ : _10844_;
  assign _10847_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [9] : \MSYNC_1r1w.synth.nz.mem[572] [9];
  assign _10848_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [9] : \MSYNC_1r1w.synth.nz.mem[574] [9];
  assign _10849_ = \bapg_rd.w_ptr_r [1] ? _10848_ : _10847_;
  assign _10850_ = \bapg_rd.w_ptr_r [2] ? _10849_ : _10846_;
  assign _10851_ = \bapg_rd.w_ptr_r [3] ? _10850_ : _10843_;
  assign _10852_ = \bapg_rd.w_ptr_r [4] ? _10851_ : _10836_;
  assign _10853_ = \bapg_rd.w_ptr_r [5] ? _10852_ : _10821_;
  assign _10854_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [9] : \MSYNC_1r1w.synth.nz.mem[576] [9];
  assign _10855_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [9] : \MSYNC_1r1w.synth.nz.mem[578] [9];
  assign _10856_ = \bapg_rd.w_ptr_r [1] ? _10855_ : _10854_;
  assign _10857_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [9] : \MSYNC_1r1w.synth.nz.mem[580] [9];
  assign _10858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [9] : \MSYNC_1r1w.synth.nz.mem[582] [9];
  assign _10859_ = \bapg_rd.w_ptr_r [1] ? _10858_ : _10857_;
  assign _10860_ = \bapg_rd.w_ptr_r [2] ? _10859_ : _10856_;
  assign _10861_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [9] : \MSYNC_1r1w.synth.nz.mem[584] [9];
  assign _10862_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [9] : \MSYNC_1r1w.synth.nz.mem[586] [9];
  assign _10863_ = \bapg_rd.w_ptr_r [1] ? _10862_ : _10861_;
  assign _10864_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [9] : \MSYNC_1r1w.synth.nz.mem[588] [9];
  assign _10865_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [9] : \MSYNC_1r1w.synth.nz.mem[590] [9];
  assign _10866_ = \bapg_rd.w_ptr_r [1] ? _10865_ : _10864_;
  assign _10867_ = \bapg_rd.w_ptr_r [2] ? _10866_ : _10863_;
  assign _10868_ = \bapg_rd.w_ptr_r [3] ? _10867_ : _10860_;
  assign _10869_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [9] : \MSYNC_1r1w.synth.nz.mem[592] [9];
  assign _10870_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [9] : \MSYNC_1r1w.synth.nz.mem[594] [9];
  assign _10871_ = \bapg_rd.w_ptr_r [1] ? _10870_ : _10869_;
  assign _10872_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [9] : \MSYNC_1r1w.synth.nz.mem[596] [9];
  assign _10873_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [9] : \MSYNC_1r1w.synth.nz.mem[598] [9];
  assign _10874_ = \bapg_rd.w_ptr_r [1] ? _10873_ : _10872_;
  assign _10875_ = \bapg_rd.w_ptr_r [2] ? _10874_ : _10871_;
  assign _10876_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [9] : \MSYNC_1r1w.synth.nz.mem[600] [9];
  assign _10877_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [9] : \MSYNC_1r1w.synth.nz.mem[602] [9];
  assign _10878_ = \bapg_rd.w_ptr_r [1] ? _10877_ : _10876_;
  assign _10879_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [9] : \MSYNC_1r1w.synth.nz.mem[604] [9];
  assign _10880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [9] : \MSYNC_1r1w.synth.nz.mem[606] [9];
  assign _10881_ = \bapg_rd.w_ptr_r [1] ? _10880_ : _10879_;
  assign _10882_ = \bapg_rd.w_ptr_r [2] ? _10881_ : _10878_;
  assign _10883_ = \bapg_rd.w_ptr_r [3] ? _10882_ : _10875_;
  assign _10884_ = \bapg_rd.w_ptr_r [4] ? _10883_ : _10868_;
  assign _10885_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [9] : \MSYNC_1r1w.synth.nz.mem[608] [9];
  assign _10886_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [9] : \MSYNC_1r1w.synth.nz.mem[610] [9];
  assign _10887_ = \bapg_rd.w_ptr_r [1] ? _10886_ : _10885_;
  assign _10888_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [9] : \MSYNC_1r1w.synth.nz.mem[612] [9];
  assign _10889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [9] : \MSYNC_1r1w.synth.nz.mem[614] [9];
  assign _10890_ = \bapg_rd.w_ptr_r [1] ? _10889_ : _10888_;
  assign _10891_ = \bapg_rd.w_ptr_r [2] ? _10890_ : _10887_;
  assign _10892_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [9] : \MSYNC_1r1w.synth.nz.mem[616] [9];
  assign _10893_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [9] : \MSYNC_1r1w.synth.nz.mem[618] [9];
  assign _10894_ = \bapg_rd.w_ptr_r [1] ? _10893_ : _10892_;
  assign _10895_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [9] : \MSYNC_1r1w.synth.nz.mem[620] [9];
  assign _10896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [9] : \MSYNC_1r1w.synth.nz.mem[622] [9];
  assign _10897_ = \bapg_rd.w_ptr_r [1] ? _10896_ : _10895_;
  assign _10898_ = \bapg_rd.w_ptr_r [2] ? _10897_ : _10894_;
  assign _10899_ = \bapg_rd.w_ptr_r [3] ? _10898_ : _10891_;
  assign _10900_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [9] : \MSYNC_1r1w.synth.nz.mem[624] [9];
  assign _10901_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [9] : \MSYNC_1r1w.synth.nz.mem[626] [9];
  assign _10902_ = \bapg_rd.w_ptr_r [1] ? _10901_ : _10900_;
  assign _10903_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [9] : \MSYNC_1r1w.synth.nz.mem[628] [9];
  assign _10904_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [9] : \MSYNC_1r1w.synth.nz.mem[630] [9];
  assign _10905_ = \bapg_rd.w_ptr_r [1] ? _10904_ : _10903_;
  assign _10906_ = \bapg_rd.w_ptr_r [2] ? _10905_ : _10902_;
  assign _10907_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [9] : \MSYNC_1r1w.synth.nz.mem[632] [9];
  assign _10908_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [9] : \MSYNC_1r1w.synth.nz.mem[634] [9];
  assign _10909_ = \bapg_rd.w_ptr_r [1] ? _10908_ : _10907_;
  assign _10910_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [9] : \MSYNC_1r1w.synth.nz.mem[636] [9];
  assign _10911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [9] : \MSYNC_1r1w.synth.nz.mem[638] [9];
  assign _10912_ = \bapg_rd.w_ptr_r [1] ? _10911_ : _10910_;
  assign _10913_ = \bapg_rd.w_ptr_r [2] ? _10912_ : _10909_;
  assign _10914_ = \bapg_rd.w_ptr_r [3] ? _10913_ : _10906_;
  assign _10915_ = \bapg_rd.w_ptr_r [4] ? _10914_ : _10899_;
  assign _10916_ = \bapg_rd.w_ptr_r [5] ? _10915_ : _10884_;
  assign _10917_ = \bapg_rd.w_ptr_r [6] ? _10916_ : _10853_;
  assign _10918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [9] : \MSYNC_1r1w.synth.nz.mem[640] [9];
  assign _10919_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [9] : \MSYNC_1r1w.synth.nz.mem[642] [9];
  assign _10920_ = \bapg_rd.w_ptr_r [1] ? _10919_ : _10918_;
  assign _10921_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [9] : \MSYNC_1r1w.synth.nz.mem[644] [9];
  assign _10922_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [9] : \MSYNC_1r1w.synth.nz.mem[646] [9];
  assign _10923_ = \bapg_rd.w_ptr_r [1] ? _10922_ : _10921_;
  assign _10924_ = \bapg_rd.w_ptr_r [2] ? _10923_ : _10920_;
  assign _10925_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [9] : \MSYNC_1r1w.synth.nz.mem[648] [9];
  assign _10926_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [9] : \MSYNC_1r1w.synth.nz.mem[650] [9];
  assign _10927_ = \bapg_rd.w_ptr_r [1] ? _10926_ : _10925_;
  assign _10928_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [9] : \MSYNC_1r1w.synth.nz.mem[652] [9];
  assign _10929_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [9] : \MSYNC_1r1w.synth.nz.mem[654] [9];
  assign _10930_ = \bapg_rd.w_ptr_r [1] ? _10929_ : _10928_;
  assign _10931_ = \bapg_rd.w_ptr_r [2] ? _10930_ : _10927_;
  assign _10932_ = \bapg_rd.w_ptr_r [3] ? _10931_ : _10924_;
  assign _10933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [9] : \MSYNC_1r1w.synth.nz.mem[656] [9];
  assign _10934_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [9] : \MSYNC_1r1w.synth.nz.mem[658] [9];
  assign _10935_ = \bapg_rd.w_ptr_r [1] ? _10934_ : _10933_;
  assign _10936_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [9] : \MSYNC_1r1w.synth.nz.mem[660] [9];
  assign _10937_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [9] : \MSYNC_1r1w.synth.nz.mem[662] [9];
  assign _10938_ = \bapg_rd.w_ptr_r [1] ? _10937_ : _10936_;
  assign _10939_ = \bapg_rd.w_ptr_r [2] ? _10938_ : _10935_;
  assign _10940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [9] : \MSYNC_1r1w.synth.nz.mem[664] [9];
  assign _10941_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [9] : \MSYNC_1r1w.synth.nz.mem[666] [9];
  assign _10942_ = \bapg_rd.w_ptr_r [1] ? _10941_ : _10940_;
  assign _10943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [9] : \MSYNC_1r1w.synth.nz.mem[668] [9];
  assign _10944_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [9] : \MSYNC_1r1w.synth.nz.mem[670] [9];
  assign _10945_ = \bapg_rd.w_ptr_r [1] ? _10944_ : _10943_;
  assign _10946_ = \bapg_rd.w_ptr_r [2] ? _10945_ : _10942_;
  assign _10947_ = \bapg_rd.w_ptr_r [3] ? _10946_ : _10939_;
  assign _10948_ = \bapg_rd.w_ptr_r [4] ? _10947_ : _10932_;
  assign _10949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [9] : \MSYNC_1r1w.synth.nz.mem[672] [9];
  assign _10950_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [9] : \MSYNC_1r1w.synth.nz.mem[674] [9];
  assign _10951_ = \bapg_rd.w_ptr_r [1] ? _10950_ : _10949_;
  assign _10952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [9] : \MSYNC_1r1w.synth.nz.mem[676] [9];
  assign _10953_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [9] : \MSYNC_1r1w.synth.nz.mem[678] [9];
  assign _10954_ = \bapg_rd.w_ptr_r [1] ? _10953_ : _10952_;
  assign _10955_ = \bapg_rd.w_ptr_r [2] ? _10954_ : _10951_;
  assign _10956_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [9] : \MSYNC_1r1w.synth.nz.mem[680] [9];
  assign _10957_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [9] : \MSYNC_1r1w.synth.nz.mem[682] [9];
  assign _10958_ = \bapg_rd.w_ptr_r [1] ? _10957_ : _10956_;
  assign _10959_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [9] : \MSYNC_1r1w.synth.nz.mem[684] [9];
  assign _10960_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [9] : \MSYNC_1r1w.synth.nz.mem[686] [9];
  assign _10961_ = \bapg_rd.w_ptr_r [1] ? _10960_ : _10959_;
  assign _10962_ = \bapg_rd.w_ptr_r [2] ? _10961_ : _10958_;
  assign _10963_ = \bapg_rd.w_ptr_r [3] ? _10962_ : _10955_;
  assign _10964_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [9] : \MSYNC_1r1w.synth.nz.mem[688] [9];
  assign _10965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [9] : \MSYNC_1r1w.synth.nz.mem[690] [9];
  assign _10966_ = \bapg_rd.w_ptr_r [1] ? _10965_ : _10964_;
  assign _10967_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [9] : \MSYNC_1r1w.synth.nz.mem[692] [9];
  assign _10968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [9] : \MSYNC_1r1w.synth.nz.mem[694] [9];
  assign _10969_ = \bapg_rd.w_ptr_r [1] ? _10968_ : _10967_;
  assign _10970_ = \bapg_rd.w_ptr_r [2] ? _10969_ : _10966_;
  assign _10971_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [9] : \MSYNC_1r1w.synth.nz.mem[696] [9];
  assign _10972_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [9] : \MSYNC_1r1w.synth.nz.mem[698] [9];
  assign _10973_ = \bapg_rd.w_ptr_r [1] ? _10972_ : _10971_;
  assign _10974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [9] : \MSYNC_1r1w.synth.nz.mem[700] [9];
  assign _10975_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [9] : \MSYNC_1r1w.synth.nz.mem[702] [9];
  assign _10976_ = \bapg_rd.w_ptr_r [1] ? _10975_ : _10974_;
  assign _10977_ = \bapg_rd.w_ptr_r [2] ? _10976_ : _10973_;
  assign _10978_ = \bapg_rd.w_ptr_r [3] ? _10977_ : _10970_;
  assign _10979_ = \bapg_rd.w_ptr_r [4] ? _10978_ : _10963_;
  assign _10980_ = \bapg_rd.w_ptr_r [5] ? _10979_ : _10948_;
  assign _10981_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [9] : \MSYNC_1r1w.synth.nz.mem[704] [9];
  assign _10982_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [9] : \MSYNC_1r1w.synth.nz.mem[706] [9];
  assign _10983_ = \bapg_rd.w_ptr_r [1] ? _10982_ : _10981_;
  assign _10984_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [9] : \MSYNC_1r1w.synth.nz.mem[708] [9];
  assign _10985_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [9] : \MSYNC_1r1w.synth.nz.mem[710] [9];
  assign _10986_ = \bapg_rd.w_ptr_r [1] ? _10985_ : _10984_;
  assign _10987_ = \bapg_rd.w_ptr_r [2] ? _10986_ : _10983_;
  assign _10988_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [9] : \MSYNC_1r1w.synth.nz.mem[712] [9];
  assign _10989_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [9] : \MSYNC_1r1w.synth.nz.mem[714] [9];
  assign _10990_ = \bapg_rd.w_ptr_r [1] ? _10989_ : _10988_;
  assign _10991_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [9] : \MSYNC_1r1w.synth.nz.mem[716] [9];
  assign _10992_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [9] : \MSYNC_1r1w.synth.nz.mem[718] [9];
  assign _10993_ = \bapg_rd.w_ptr_r [1] ? _10992_ : _10991_;
  assign _10994_ = \bapg_rd.w_ptr_r [2] ? _10993_ : _10990_;
  assign _10995_ = \bapg_rd.w_ptr_r [3] ? _10994_ : _10987_;
  assign _10996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [9] : \MSYNC_1r1w.synth.nz.mem[720] [9];
  assign _10997_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [9] : \MSYNC_1r1w.synth.nz.mem[722] [9];
  assign _10998_ = \bapg_rd.w_ptr_r [1] ? _10997_ : _10996_;
  assign _10999_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [9] : \MSYNC_1r1w.synth.nz.mem[724] [9];
  assign _11000_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [9] : \MSYNC_1r1w.synth.nz.mem[726] [9];
  assign _11001_ = \bapg_rd.w_ptr_r [1] ? _11000_ : _10999_;
  assign _11002_ = \bapg_rd.w_ptr_r [2] ? _11001_ : _10998_;
  assign _11003_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [9] : \MSYNC_1r1w.synth.nz.mem[728] [9];
  assign _11004_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [9] : \MSYNC_1r1w.synth.nz.mem[730] [9];
  assign _11005_ = \bapg_rd.w_ptr_r [1] ? _11004_ : _11003_;
  assign _11006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [9] : \MSYNC_1r1w.synth.nz.mem[732] [9];
  assign _11007_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [9] : \MSYNC_1r1w.synth.nz.mem[734] [9];
  assign _11008_ = \bapg_rd.w_ptr_r [1] ? _11007_ : _11006_;
  assign _11009_ = \bapg_rd.w_ptr_r [2] ? _11008_ : _11005_;
  assign _11010_ = \bapg_rd.w_ptr_r [3] ? _11009_ : _11002_;
  assign _11011_ = \bapg_rd.w_ptr_r [4] ? _11010_ : _10995_;
  assign _11012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [9] : \MSYNC_1r1w.synth.nz.mem[736] [9];
  assign _11013_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [9] : \MSYNC_1r1w.synth.nz.mem[738] [9];
  assign _11014_ = \bapg_rd.w_ptr_r [1] ? _11013_ : _11012_;
  assign _11015_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [9] : \MSYNC_1r1w.synth.nz.mem[740] [9];
  assign _11016_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [9] : \MSYNC_1r1w.synth.nz.mem[742] [9];
  assign _11017_ = \bapg_rd.w_ptr_r [1] ? _11016_ : _11015_;
  assign _11018_ = \bapg_rd.w_ptr_r [2] ? _11017_ : _11014_;
  assign _11019_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [9] : \MSYNC_1r1w.synth.nz.mem[744] [9];
  assign _11020_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [9] : \MSYNC_1r1w.synth.nz.mem[746] [9];
  assign _11021_ = \bapg_rd.w_ptr_r [1] ? _11020_ : _11019_;
  assign _11022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [9] : \MSYNC_1r1w.synth.nz.mem[748] [9];
  assign _11023_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [9] : \MSYNC_1r1w.synth.nz.mem[750] [9];
  assign _11024_ = \bapg_rd.w_ptr_r [1] ? _11023_ : _11022_;
  assign _11025_ = \bapg_rd.w_ptr_r [2] ? _11024_ : _11021_;
  assign _11026_ = \bapg_rd.w_ptr_r [3] ? _11025_ : _11018_;
  assign _11027_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [9] : \MSYNC_1r1w.synth.nz.mem[752] [9];
  assign _11028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [9] : \MSYNC_1r1w.synth.nz.mem[754] [9];
  assign _11029_ = \bapg_rd.w_ptr_r [1] ? _11028_ : _11027_;
  assign _11030_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [9] : \MSYNC_1r1w.synth.nz.mem[756] [9];
  assign _11031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [9] : \MSYNC_1r1w.synth.nz.mem[758] [9];
  assign _11032_ = \bapg_rd.w_ptr_r [1] ? _11031_ : _11030_;
  assign _11033_ = \bapg_rd.w_ptr_r [2] ? _11032_ : _11029_;
  assign _11034_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [9] : \MSYNC_1r1w.synth.nz.mem[760] [9];
  assign _11035_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [9] : \MSYNC_1r1w.synth.nz.mem[762] [9];
  assign _11036_ = \bapg_rd.w_ptr_r [1] ? _11035_ : _11034_;
  assign _11037_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [9] : \MSYNC_1r1w.synth.nz.mem[764] [9];
  assign _11038_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [9] : \MSYNC_1r1w.synth.nz.mem[766] [9];
  assign _11039_ = \bapg_rd.w_ptr_r [1] ? _11038_ : _11037_;
  assign _11040_ = \bapg_rd.w_ptr_r [2] ? _11039_ : _11036_;
  assign _11041_ = \bapg_rd.w_ptr_r [3] ? _11040_ : _11033_;
  assign _11042_ = \bapg_rd.w_ptr_r [4] ? _11041_ : _11026_;
  assign _11043_ = \bapg_rd.w_ptr_r [5] ? _11042_ : _11011_;
  assign _11044_ = \bapg_rd.w_ptr_r [6] ? _11043_ : _10980_;
  assign _11045_ = \bapg_rd.w_ptr_r [7] ? _11044_ : _10917_;
  assign _11046_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [9] : \MSYNC_1r1w.synth.nz.mem[768] [9];
  assign _11047_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [9] : \MSYNC_1r1w.synth.nz.mem[770] [9];
  assign _11048_ = \bapg_rd.w_ptr_r [1] ? _11047_ : _11046_;
  assign _11049_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [9] : \MSYNC_1r1w.synth.nz.mem[772] [9];
  assign _11050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [9] : \MSYNC_1r1w.synth.nz.mem[774] [9];
  assign _11051_ = \bapg_rd.w_ptr_r [1] ? _11050_ : _11049_;
  assign _11052_ = \bapg_rd.w_ptr_r [2] ? _11051_ : _11048_;
  assign _11053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [9] : \MSYNC_1r1w.synth.nz.mem[776] [9];
  assign _11054_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [9] : \MSYNC_1r1w.synth.nz.mem[778] [9];
  assign _11055_ = \bapg_rd.w_ptr_r [1] ? _11054_ : _11053_;
  assign _11056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [9] : \MSYNC_1r1w.synth.nz.mem[780] [9];
  assign _11057_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [9] : \MSYNC_1r1w.synth.nz.mem[782] [9];
  assign _11058_ = \bapg_rd.w_ptr_r [1] ? _11057_ : _11056_;
  assign _11059_ = \bapg_rd.w_ptr_r [2] ? _11058_ : _11055_;
  assign _11060_ = \bapg_rd.w_ptr_r [3] ? _11059_ : _11052_;
  assign _11061_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [9] : \MSYNC_1r1w.synth.nz.mem[784] [9];
  assign _11062_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [9] : \MSYNC_1r1w.synth.nz.mem[786] [9];
  assign _11063_ = \bapg_rd.w_ptr_r [1] ? _11062_ : _11061_;
  assign _11064_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [9] : \MSYNC_1r1w.synth.nz.mem[788] [9];
  assign _11065_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [9] : \MSYNC_1r1w.synth.nz.mem[790] [9];
  assign _11066_ = \bapg_rd.w_ptr_r [1] ? _11065_ : _11064_;
  assign _11067_ = \bapg_rd.w_ptr_r [2] ? _11066_ : _11063_;
  assign _11068_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [9] : \MSYNC_1r1w.synth.nz.mem[792] [9];
  assign _11069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [9] : \MSYNC_1r1w.synth.nz.mem[794] [9];
  assign _11070_ = \bapg_rd.w_ptr_r [1] ? _11069_ : _11068_;
  assign _11071_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [9] : \MSYNC_1r1w.synth.nz.mem[796] [9];
  assign _11072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [9] : \MSYNC_1r1w.synth.nz.mem[798] [9];
  assign _11073_ = \bapg_rd.w_ptr_r [1] ? _11072_ : _11071_;
  assign _11074_ = \bapg_rd.w_ptr_r [2] ? _11073_ : _11070_;
  assign _11075_ = \bapg_rd.w_ptr_r [3] ? _11074_ : _11067_;
  assign _11076_ = \bapg_rd.w_ptr_r [4] ? _11075_ : _11060_;
  assign _11077_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [9] : \MSYNC_1r1w.synth.nz.mem[800] [9];
  assign _11078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [9] : \MSYNC_1r1w.synth.nz.mem[802] [9];
  assign _11079_ = \bapg_rd.w_ptr_r [1] ? _11078_ : _11077_;
  assign _11080_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [9] : \MSYNC_1r1w.synth.nz.mem[804] [9];
  assign _11081_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [9] : \MSYNC_1r1w.synth.nz.mem[806] [9];
  assign _11082_ = \bapg_rd.w_ptr_r [1] ? _11081_ : _11080_;
  assign _11083_ = \bapg_rd.w_ptr_r [2] ? _11082_ : _11079_;
  assign _11084_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [9] : \MSYNC_1r1w.synth.nz.mem[808] [9];
  assign _11085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [9] : \MSYNC_1r1w.synth.nz.mem[810] [9];
  assign _11086_ = \bapg_rd.w_ptr_r [1] ? _11085_ : _11084_;
  assign _11087_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [9] : \MSYNC_1r1w.synth.nz.mem[812] [9];
  assign _11088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [9] : \MSYNC_1r1w.synth.nz.mem[814] [9];
  assign _11089_ = \bapg_rd.w_ptr_r [1] ? _11088_ : _11087_;
  assign _11090_ = \bapg_rd.w_ptr_r [2] ? _11089_ : _11086_;
  assign _11091_ = \bapg_rd.w_ptr_r [3] ? _11090_ : _11083_;
  assign _11092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [9] : \MSYNC_1r1w.synth.nz.mem[816] [9];
  assign _11093_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [9] : \MSYNC_1r1w.synth.nz.mem[818] [9];
  assign _11094_ = \bapg_rd.w_ptr_r [1] ? _11093_ : _11092_;
  assign _11095_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [9] : \MSYNC_1r1w.synth.nz.mem[820] [9];
  assign _11096_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [9] : \MSYNC_1r1w.synth.nz.mem[822] [9];
  assign _11097_ = \bapg_rd.w_ptr_r [1] ? _11096_ : _11095_;
  assign _11098_ = \bapg_rd.w_ptr_r [2] ? _11097_ : _11094_;
  assign _11099_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [9] : \MSYNC_1r1w.synth.nz.mem[824] [9];
  assign _11100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [9] : \MSYNC_1r1w.synth.nz.mem[826] [9];
  assign _11101_ = \bapg_rd.w_ptr_r [1] ? _11100_ : _11099_;
  assign _11102_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [9] : \MSYNC_1r1w.synth.nz.mem[828] [9];
  assign _11103_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [9] : \MSYNC_1r1w.synth.nz.mem[830] [9];
  assign _11104_ = \bapg_rd.w_ptr_r [1] ? _11103_ : _11102_;
  assign _11105_ = \bapg_rd.w_ptr_r [2] ? _11104_ : _11101_;
  assign _11106_ = \bapg_rd.w_ptr_r [3] ? _11105_ : _11098_;
  assign _11107_ = \bapg_rd.w_ptr_r [4] ? _11106_ : _11091_;
  assign _11108_ = \bapg_rd.w_ptr_r [5] ? _11107_ : _11076_;
  assign _11109_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [9] : \MSYNC_1r1w.synth.nz.mem[832] [9];
  assign _11110_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [9] : \MSYNC_1r1w.synth.nz.mem[834] [9];
  assign _11111_ = \bapg_rd.w_ptr_r [1] ? _11110_ : _11109_;
  assign _11112_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [9] : \MSYNC_1r1w.synth.nz.mem[836] [9];
  assign _11113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [9] : \MSYNC_1r1w.synth.nz.mem[838] [9];
  assign _11114_ = \bapg_rd.w_ptr_r [1] ? _11113_ : _11112_;
  assign _11115_ = \bapg_rd.w_ptr_r [2] ? _11114_ : _11111_;
  assign _11116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [9] : \MSYNC_1r1w.synth.nz.mem[840] [9];
  assign _11117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [9] : \MSYNC_1r1w.synth.nz.mem[842] [9];
  assign _11118_ = \bapg_rd.w_ptr_r [1] ? _11117_ : _11116_;
  assign _11119_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [9] : \MSYNC_1r1w.synth.nz.mem[844] [9];
  assign _11120_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [9] : \MSYNC_1r1w.synth.nz.mem[846] [9];
  assign _11121_ = \bapg_rd.w_ptr_r [1] ? _11120_ : _11119_;
  assign _11122_ = \bapg_rd.w_ptr_r [2] ? _11121_ : _11118_;
  assign _11123_ = \bapg_rd.w_ptr_r [3] ? _11122_ : _11115_;
  assign _11124_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [9] : \MSYNC_1r1w.synth.nz.mem[848] [9];
  assign _11125_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [9] : \MSYNC_1r1w.synth.nz.mem[850] [9];
  assign _11126_ = \bapg_rd.w_ptr_r [1] ? _11125_ : _11124_;
  assign _11127_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [9] : \MSYNC_1r1w.synth.nz.mem[852] [9];
  assign _11128_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [9] : \MSYNC_1r1w.synth.nz.mem[854] [9];
  assign _11129_ = \bapg_rd.w_ptr_r [1] ? _11128_ : _11127_;
  assign _11130_ = \bapg_rd.w_ptr_r [2] ? _11129_ : _11126_;
  assign _11131_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [9] : \MSYNC_1r1w.synth.nz.mem[856] [9];
  assign _11132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [9] : \MSYNC_1r1w.synth.nz.mem[858] [9];
  assign _11133_ = \bapg_rd.w_ptr_r [1] ? _11132_ : _11131_;
  assign _11134_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [9] : \MSYNC_1r1w.synth.nz.mem[860] [9];
  assign _11135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [9] : \MSYNC_1r1w.synth.nz.mem[862] [9];
  assign _11136_ = \bapg_rd.w_ptr_r [1] ? _11135_ : _11134_;
  assign _11137_ = \bapg_rd.w_ptr_r [2] ? _11136_ : _11133_;
  assign _11138_ = \bapg_rd.w_ptr_r [3] ? _11137_ : _11130_;
  assign _11139_ = \bapg_rd.w_ptr_r [4] ? _11138_ : _11123_;
  assign _11140_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [9] : \MSYNC_1r1w.synth.nz.mem[864] [9];
  assign _11141_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [9] : \MSYNC_1r1w.synth.nz.mem[866] [9];
  assign _11142_ = \bapg_rd.w_ptr_r [1] ? _11141_ : _11140_;
  assign _11143_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [9] : \MSYNC_1r1w.synth.nz.mem[868] [9];
  assign _11144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [9] : \MSYNC_1r1w.synth.nz.mem[870] [9];
  assign _11145_ = \bapg_rd.w_ptr_r [1] ? _11144_ : _11143_;
  assign _11146_ = \bapg_rd.w_ptr_r [2] ? _11145_ : _11142_;
  assign _11147_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [9] : \MSYNC_1r1w.synth.nz.mem[872] [9];
  assign _11148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [9] : \MSYNC_1r1w.synth.nz.mem[874] [9];
  assign _11149_ = \bapg_rd.w_ptr_r [1] ? _11148_ : _11147_;
  assign _11150_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [9] : \MSYNC_1r1w.synth.nz.mem[876] [9];
  assign _11151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [9] : \MSYNC_1r1w.synth.nz.mem[878] [9];
  assign _11152_ = \bapg_rd.w_ptr_r [1] ? _11151_ : _11150_;
  assign _11153_ = \bapg_rd.w_ptr_r [2] ? _11152_ : _11149_;
  assign _11154_ = \bapg_rd.w_ptr_r [3] ? _11153_ : _11146_;
  assign _11155_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [9] : \MSYNC_1r1w.synth.nz.mem[880] [9];
  assign _11156_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [9] : \MSYNC_1r1w.synth.nz.mem[882] [9];
  assign _11157_ = \bapg_rd.w_ptr_r [1] ? _11156_ : _11155_;
  assign _11158_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [9] : \MSYNC_1r1w.synth.nz.mem[884] [9];
  assign _11159_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [9] : \MSYNC_1r1w.synth.nz.mem[886] [9];
  assign _11160_ = \bapg_rd.w_ptr_r [1] ? _11159_ : _11158_;
  assign _11161_ = \bapg_rd.w_ptr_r [2] ? _11160_ : _11157_;
  assign _11162_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [9] : \MSYNC_1r1w.synth.nz.mem[888] [9];
  assign _11163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [9] : \MSYNC_1r1w.synth.nz.mem[890] [9];
  assign _11164_ = \bapg_rd.w_ptr_r [1] ? _11163_ : _11162_;
  assign _11165_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [9] : \MSYNC_1r1w.synth.nz.mem[892] [9];
  assign _11166_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [9] : \MSYNC_1r1w.synth.nz.mem[894] [9];
  assign _11167_ = \bapg_rd.w_ptr_r [1] ? _11166_ : _11165_;
  assign _11168_ = \bapg_rd.w_ptr_r [2] ? _11167_ : _11164_;
  assign _11169_ = \bapg_rd.w_ptr_r [3] ? _11168_ : _11161_;
  assign _11170_ = \bapg_rd.w_ptr_r [4] ? _11169_ : _11154_;
  assign _11171_ = \bapg_rd.w_ptr_r [5] ? _11170_ : _11139_;
  assign _11172_ = \bapg_rd.w_ptr_r [6] ? _11171_ : _11108_;
  assign _11173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [9] : \MSYNC_1r1w.synth.nz.mem[896] [9];
  assign _11174_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [9] : \MSYNC_1r1w.synth.nz.mem[898] [9];
  assign _11175_ = \bapg_rd.w_ptr_r [1] ? _11174_ : _11173_;
  assign _11176_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [9] : \MSYNC_1r1w.synth.nz.mem[900] [9];
  assign _11177_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [9] : \MSYNC_1r1w.synth.nz.mem[902] [9];
  assign _11178_ = \bapg_rd.w_ptr_r [1] ? _11177_ : _11176_;
  assign _11179_ = \bapg_rd.w_ptr_r [2] ? _11178_ : _11175_;
  assign _11180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [9] : \MSYNC_1r1w.synth.nz.mem[904] [9];
  assign _11181_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [9] : \MSYNC_1r1w.synth.nz.mem[906] [9];
  assign _11182_ = \bapg_rd.w_ptr_r [1] ? _11181_ : _11180_;
  assign _11183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [9] : \MSYNC_1r1w.synth.nz.mem[908] [9];
  assign _11184_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [9] : \MSYNC_1r1w.synth.nz.mem[910] [9];
  assign _11185_ = \bapg_rd.w_ptr_r [1] ? _11184_ : _11183_;
  assign _11186_ = \bapg_rd.w_ptr_r [2] ? _11185_ : _11182_;
  assign _11187_ = \bapg_rd.w_ptr_r [3] ? _11186_ : _11179_;
  assign _11188_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [9] : \MSYNC_1r1w.synth.nz.mem[912] [9];
  assign _11189_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [9] : \MSYNC_1r1w.synth.nz.mem[914] [9];
  assign _11190_ = \bapg_rd.w_ptr_r [1] ? _11189_ : _11188_;
  assign _11191_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [9] : \MSYNC_1r1w.synth.nz.mem[916] [9];
  assign _11192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [9] : \MSYNC_1r1w.synth.nz.mem[918] [9];
  assign _11193_ = \bapg_rd.w_ptr_r [1] ? _11192_ : _11191_;
  assign _11194_ = \bapg_rd.w_ptr_r [2] ? _11193_ : _11190_;
  assign _11195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [9] : \MSYNC_1r1w.synth.nz.mem[920] [9];
  assign _11196_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [9] : \MSYNC_1r1w.synth.nz.mem[922] [9];
  assign _11197_ = \bapg_rd.w_ptr_r [1] ? _11196_ : _11195_;
  assign _11198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [9] : \MSYNC_1r1w.synth.nz.mem[924] [9];
  assign _11199_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [9] : \MSYNC_1r1w.synth.nz.mem[926] [9];
  assign _11200_ = \bapg_rd.w_ptr_r [1] ? _11199_ : _11198_;
  assign _11201_ = \bapg_rd.w_ptr_r [2] ? _11200_ : _11197_;
  assign _11202_ = \bapg_rd.w_ptr_r [3] ? _11201_ : _11194_;
  assign _11203_ = \bapg_rd.w_ptr_r [4] ? _11202_ : _11187_;
  assign _11204_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [9] : \MSYNC_1r1w.synth.nz.mem[928] [9];
  assign _11205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [9] : \MSYNC_1r1w.synth.nz.mem[930] [9];
  assign _11206_ = \bapg_rd.w_ptr_r [1] ? _11205_ : _11204_;
  assign _11207_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [9] : \MSYNC_1r1w.synth.nz.mem[932] [9];
  assign _11208_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [9] : \MSYNC_1r1w.synth.nz.mem[934] [9];
  assign _11209_ = \bapg_rd.w_ptr_r [1] ? _11208_ : _11207_;
  assign _11210_ = \bapg_rd.w_ptr_r [2] ? _11209_ : _11206_;
  assign _11211_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [9] : \MSYNC_1r1w.synth.nz.mem[936] [9];
  assign _11212_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [9] : \MSYNC_1r1w.synth.nz.mem[938] [9];
  assign _11213_ = \bapg_rd.w_ptr_r [1] ? _11212_ : _11211_;
  assign _11214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [9] : \MSYNC_1r1w.synth.nz.mem[940] [9];
  assign _11215_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [9] : \MSYNC_1r1w.synth.nz.mem[942] [9];
  assign _11216_ = \bapg_rd.w_ptr_r [1] ? _11215_ : _11214_;
  assign _11217_ = \bapg_rd.w_ptr_r [2] ? _11216_ : _11213_;
  assign _11218_ = \bapg_rd.w_ptr_r [3] ? _11217_ : _11210_;
  assign _11219_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [9] : \MSYNC_1r1w.synth.nz.mem[944] [9];
  assign _11220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [9] : \MSYNC_1r1w.synth.nz.mem[946] [9];
  assign _11221_ = \bapg_rd.w_ptr_r [1] ? _11220_ : _11219_;
  assign _11222_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [9] : \MSYNC_1r1w.synth.nz.mem[948] [9];
  assign _11223_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [9] : \MSYNC_1r1w.synth.nz.mem[950] [9];
  assign _11224_ = \bapg_rd.w_ptr_r [1] ? _11223_ : _11222_;
  assign _11225_ = \bapg_rd.w_ptr_r [2] ? _11224_ : _11221_;
  assign _11226_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [9] : \MSYNC_1r1w.synth.nz.mem[952] [9];
  assign _11227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [9] : \MSYNC_1r1w.synth.nz.mem[954] [9];
  assign _11228_ = \bapg_rd.w_ptr_r [1] ? _11227_ : _11226_;
  assign _11229_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [9] : \MSYNC_1r1w.synth.nz.mem[956] [9];
  assign _11230_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [9] : \MSYNC_1r1w.synth.nz.mem[958] [9];
  assign _11231_ = \bapg_rd.w_ptr_r [1] ? _11230_ : _11229_;
  assign _11232_ = \bapg_rd.w_ptr_r [2] ? _11231_ : _11228_;
  assign _11233_ = \bapg_rd.w_ptr_r [3] ? _11232_ : _11225_;
  assign _11234_ = \bapg_rd.w_ptr_r [4] ? _11233_ : _11218_;
  assign _11235_ = \bapg_rd.w_ptr_r [5] ? _11234_ : _11203_;
  assign _11236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [9] : \MSYNC_1r1w.synth.nz.mem[960] [9];
  assign _11237_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [9] : \MSYNC_1r1w.synth.nz.mem[962] [9];
  assign _11238_ = \bapg_rd.w_ptr_r [1] ? _11237_ : _11236_;
  assign _11239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [9] : \MSYNC_1r1w.synth.nz.mem[964] [9];
  assign _11240_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [9] : \MSYNC_1r1w.synth.nz.mem[966] [9];
  assign _11241_ = \bapg_rd.w_ptr_r [1] ? _11240_ : _11239_;
  assign _11242_ = \bapg_rd.w_ptr_r [2] ? _11241_ : _11238_;
  assign _11243_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [9] : \MSYNC_1r1w.synth.nz.mem[968] [9];
  assign _11244_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [9] : \MSYNC_1r1w.synth.nz.mem[970] [9];
  assign _11245_ = \bapg_rd.w_ptr_r [1] ? _11244_ : _11243_;
  assign _11246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [9] : \MSYNC_1r1w.synth.nz.mem[972] [9];
  assign _11247_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [9] : \MSYNC_1r1w.synth.nz.mem[974] [9];
  assign _11248_ = \bapg_rd.w_ptr_r [1] ? _11247_ : _11246_;
  assign _11249_ = \bapg_rd.w_ptr_r [2] ? _11248_ : _11245_;
  assign _11250_ = \bapg_rd.w_ptr_r [3] ? _11249_ : _11242_;
  assign _11251_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [9] : \MSYNC_1r1w.synth.nz.mem[976] [9];
  assign _11252_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [9] : \MSYNC_1r1w.synth.nz.mem[978] [9];
  assign _11253_ = \bapg_rd.w_ptr_r [1] ? _11252_ : _11251_;
  assign _11254_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [9] : \MSYNC_1r1w.synth.nz.mem[980] [9];
  assign _11255_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [9] : \MSYNC_1r1w.synth.nz.mem[982] [9];
  assign _11256_ = \bapg_rd.w_ptr_r [1] ? _11255_ : _11254_;
  assign _11257_ = \bapg_rd.w_ptr_r [2] ? _11256_ : _11253_;
  assign _11258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [9] : \MSYNC_1r1w.synth.nz.mem[984] [9];
  assign _11259_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [9] : \MSYNC_1r1w.synth.nz.mem[986] [9];
  assign _11260_ = \bapg_rd.w_ptr_r [1] ? _11259_ : _11258_;
  assign _11261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [9] : \MSYNC_1r1w.synth.nz.mem[988] [9];
  assign _11262_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [9] : \MSYNC_1r1w.synth.nz.mem[990] [9];
  assign _11263_ = \bapg_rd.w_ptr_r [1] ? _11262_ : _11261_;
  assign _11264_ = \bapg_rd.w_ptr_r [2] ? _11263_ : _11260_;
  assign _11265_ = \bapg_rd.w_ptr_r [3] ? _11264_ : _11257_;
  assign _11266_ = \bapg_rd.w_ptr_r [4] ? _11265_ : _11250_;
  assign _11267_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [9] : \MSYNC_1r1w.synth.nz.mem[992] [9];
  assign _11268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [9] : \MSYNC_1r1w.synth.nz.mem[994] [9];
  assign _11269_ = \bapg_rd.w_ptr_r [1] ? _11268_ : _11267_;
  assign _11270_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [9] : \MSYNC_1r1w.synth.nz.mem[996] [9];
  assign _11271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [9] : \MSYNC_1r1w.synth.nz.mem[998] [9];
  assign _11272_ = \bapg_rd.w_ptr_r [1] ? _11271_ : _11270_;
  assign _11273_ = \bapg_rd.w_ptr_r [2] ? _11272_ : _11269_;
  assign _11274_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [9] : \MSYNC_1r1w.synth.nz.mem[1000] [9];
  assign _11275_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [9] : \MSYNC_1r1w.synth.nz.mem[1002] [9];
  assign _11276_ = \bapg_rd.w_ptr_r [1] ? _11275_ : _11274_;
  assign _11277_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [9] : \MSYNC_1r1w.synth.nz.mem[1004] [9];
  assign _11278_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [9] : \MSYNC_1r1w.synth.nz.mem[1006] [9];
  assign _11279_ = \bapg_rd.w_ptr_r [1] ? _11278_ : _11277_;
  assign _11280_ = \bapg_rd.w_ptr_r [2] ? _11279_ : _11276_;
  assign _11281_ = \bapg_rd.w_ptr_r [3] ? _11280_ : _11273_;
  assign _11282_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [9] : \MSYNC_1r1w.synth.nz.mem[1008] [9];
  assign _11283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [9] : \MSYNC_1r1w.synth.nz.mem[1010] [9];
  assign _11284_ = \bapg_rd.w_ptr_r [1] ? _11283_ : _11282_;
  assign _11285_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [9] : \MSYNC_1r1w.synth.nz.mem[1012] [9];
  assign _11286_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [9] : \MSYNC_1r1w.synth.nz.mem[1014] [9];
  assign _11287_ = \bapg_rd.w_ptr_r [1] ? _11286_ : _11285_;
  assign _11288_ = \bapg_rd.w_ptr_r [2] ? _11287_ : _11284_;
  assign _11289_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [9] : \MSYNC_1r1w.synth.nz.mem[1016] [9];
  assign _11290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [9] : \MSYNC_1r1w.synth.nz.mem[1018] [9];
  assign _11291_ = \bapg_rd.w_ptr_r [1] ? _11290_ : _11289_;
  assign _11292_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [9] : \MSYNC_1r1w.synth.nz.mem[1020] [9];
  assign _11293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [9] : \MSYNC_1r1w.synth.nz.mem[1022] [9];
  assign _11294_ = \bapg_rd.w_ptr_r [1] ? _11293_ : _11292_;
  assign _11295_ = \bapg_rd.w_ptr_r [2] ? _11294_ : _11291_;
  assign _11296_ = \bapg_rd.w_ptr_r [3] ? _11295_ : _11288_;
  assign _11297_ = \bapg_rd.w_ptr_r [4] ? _11296_ : _11281_;
  assign _11298_ = \bapg_rd.w_ptr_r [5] ? _11297_ : _11266_;
  assign _11299_ = \bapg_rd.w_ptr_r [6] ? _11298_ : _11235_;
  assign _11300_ = \bapg_rd.w_ptr_r [7] ? _11299_ : _11172_;
  assign _11301_ = \bapg_rd.w_ptr_r [8] ? _11300_ : _11045_;
  assign r_data_o[9] = \bapg_rd.w_ptr_r [9] ? _11301_ : _10790_;
  assign _11302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [10] : \MSYNC_1r1w.synth.nz.mem[0] [10];
  assign _11303_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [10] : \MSYNC_1r1w.synth.nz.mem[2] [10];
  assign _11304_ = \bapg_rd.w_ptr_r [1] ? _11303_ : _11302_;
  assign _11305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [10] : \MSYNC_1r1w.synth.nz.mem[4] [10];
  assign _11306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [10] : \MSYNC_1r1w.synth.nz.mem[6] [10];
  assign _11307_ = \bapg_rd.w_ptr_r [1] ? _11306_ : _11305_;
  assign _11308_ = \bapg_rd.w_ptr_r [2] ? _11307_ : _11304_;
  assign _11309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [10] : \MSYNC_1r1w.synth.nz.mem[8] [10];
  assign _11310_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [10] : \MSYNC_1r1w.synth.nz.mem[10] [10];
  assign _11311_ = \bapg_rd.w_ptr_r [1] ? _11310_ : _11309_;
  assign _11312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [10] : \MSYNC_1r1w.synth.nz.mem[12] [10];
  assign _11313_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [10] : \MSYNC_1r1w.synth.nz.mem[14] [10];
  assign _11314_ = \bapg_rd.w_ptr_r [1] ? _11313_ : _11312_;
  assign _11315_ = \bapg_rd.w_ptr_r [2] ? _11314_ : _11311_;
  assign _11316_ = \bapg_rd.w_ptr_r [3] ? _11315_ : _11308_;
  assign _11317_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [10] : \MSYNC_1r1w.synth.nz.mem[16] [10];
  assign _11318_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [10] : \MSYNC_1r1w.synth.nz.mem[18] [10];
  assign _11319_ = \bapg_rd.w_ptr_r [1] ? _11318_ : _11317_;
  assign _11320_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [10] : \MSYNC_1r1w.synth.nz.mem[20] [10];
  assign _11321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [10] : \MSYNC_1r1w.synth.nz.mem[22] [10];
  assign _11322_ = \bapg_rd.w_ptr_r [1] ? _11321_ : _11320_;
  assign _11323_ = \bapg_rd.w_ptr_r [2] ? _11322_ : _11319_;
  assign _11324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [10] : \MSYNC_1r1w.synth.nz.mem[24] [10];
  assign _11325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [10] : \MSYNC_1r1w.synth.nz.mem[26] [10];
  assign _11326_ = \bapg_rd.w_ptr_r [1] ? _11325_ : _11324_;
  assign _11327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [10] : \MSYNC_1r1w.synth.nz.mem[28] [10];
  assign _11328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [10] : \MSYNC_1r1w.synth.nz.mem[30] [10];
  assign _11329_ = \bapg_rd.w_ptr_r [1] ? _11328_ : _11327_;
  assign _11330_ = \bapg_rd.w_ptr_r [2] ? _11329_ : _11326_;
  assign _11331_ = \bapg_rd.w_ptr_r [3] ? _11330_ : _11323_;
  assign _11332_ = \bapg_rd.w_ptr_r [4] ? _11331_ : _11316_;
  assign _11333_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [10] : \MSYNC_1r1w.synth.nz.mem[32] [10];
  assign _11334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [10] : \MSYNC_1r1w.synth.nz.mem[34] [10];
  assign _11335_ = \bapg_rd.w_ptr_r [1] ? _11334_ : _11333_;
  assign _11336_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [10] : \MSYNC_1r1w.synth.nz.mem[36] [10];
  assign _11337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [10] : \MSYNC_1r1w.synth.nz.mem[38] [10];
  assign _11338_ = \bapg_rd.w_ptr_r [1] ? _11337_ : _11336_;
  assign _11339_ = \bapg_rd.w_ptr_r [2] ? _11338_ : _11335_;
  assign _11340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [10] : \MSYNC_1r1w.synth.nz.mem[40] [10];
  assign _11341_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [10] : \MSYNC_1r1w.synth.nz.mem[42] [10];
  assign _11342_ = \bapg_rd.w_ptr_r [1] ? _11341_ : _11340_;
  assign _11343_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [10] : \MSYNC_1r1w.synth.nz.mem[44] [10];
  assign _11344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [10] : \MSYNC_1r1w.synth.nz.mem[46] [10];
  assign _11345_ = \bapg_rd.w_ptr_r [1] ? _11344_ : _11343_;
  assign _11346_ = \bapg_rd.w_ptr_r [2] ? _11345_ : _11342_;
  assign _11347_ = \bapg_rd.w_ptr_r [3] ? _11346_ : _11339_;
  assign _11348_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [10] : \MSYNC_1r1w.synth.nz.mem[48] [10];
  assign _11349_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [10] : \MSYNC_1r1w.synth.nz.mem[50] [10];
  assign _11350_ = \bapg_rd.w_ptr_r [1] ? _11349_ : _11348_;
  assign _11351_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [10] : \MSYNC_1r1w.synth.nz.mem[52] [10];
  assign _11352_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [10] : \MSYNC_1r1w.synth.nz.mem[54] [10];
  assign _11353_ = \bapg_rd.w_ptr_r [1] ? _11352_ : _11351_;
  assign _11354_ = \bapg_rd.w_ptr_r [2] ? _11353_ : _11350_;
  assign _11355_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [10] : \MSYNC_1r1w.synth.nz.mem[56] [10];
  assign _11356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [10] : \MSYNC_1r1w.synth.nz.mem[58] [10];
  assign _11357_ = \bapg_rd.w_ptr_r [1] ? _11356_ : _11355_;
  assign _11358_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [10] : \MSYNC_1r1w.synth.nz.mem[60] [10];
  assign _11359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [10] : \MSYNC_1r1w.synth.nz.mem[62] [10];
  assign _11360_ = \bapg_rd.w_ptr_r [1] ? _11359_ : _11358_;
  assign _11361_ = \bapg_rd.w_ptr_r [2] ? _11360_ : _11357_;
  assign _11362_ = \bapg_rd.w_ptr_r [3] ? _11361_ : _11354_;
  assign _11363_ = \bapg_rd.w_ptr_r [4] ? _11362_ : _11347_;
  assign _11364_ = \bapg_rd.w_ptr_r [5] ? _11363_ : _11332_;
  assign _11365_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [10] : \MSYNC_1r1w.synth.nz.mem[64] [10];
  assign _11366_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [10] : \MSYNC_1r1w.synth.nz.mem[66] [10];
  assign _11367_ = \bapg_rd.w_ptr_r [1] ? _11366_ : _11365_;
  assign _11368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [10] : \MSYNC_1r1w.synth.nz.mem[68] [10];
  assign _11369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [10] : \MSYNC_1r1w.synth.nz.mem[70] [10];
  assign _11370_ = \bapg_rd.w_ptr_r [1] ? _11369_ : _11368_;
  assign _11371_ = \bapg_rd.w_ptr_r [2] ? _11370_ : _11367_;
  assign _11372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [10] : \MSYNC_1r1w.synth.nz.mem[72] [10];
  assign _11373_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [10] : \MSYNC_1r1w.synth.nz.mem[74] [10];
  assign _11374_ = \bapg_rd.w_ptr_r [1] ? _11373_ : _11372_;
  assign _11375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [10] : \MSYNC_1r1w.synth.nz.mem[76] [10];
  assign _11376_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [10] : \MSYNC_1r1w.synth.nz.mem[78] [10];
  assign _11377_ = \bapg_rd.w_ptr_r [1] ? _11376_ : _11375_;
  assign _11378_ = \bapg_rd.w_ptr_r [2] ? _11377_ : _11374_;
  assign _11379_ = \bapg_rd.w_ptr_r [3] ? _11378_ : _11371_;
  assign _11380_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [10] : \MSYNC_1r1w.synth.nz.mem[80] [10];
  assign _11381_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [10] : \MSYNC_1r1w.synth.nz.mem[82] [10];
  assign _11382_ = \bapg_rd.w_ptr_r [1] ? _11381_ : _11380_;
  assign _11383_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [10] : \MSYNC_1r1w.synth.nz.mem[84] [10];
  assign _11384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [10] : \MSYNC_1r1w.synth.nz.mem[86] [10];
  assign _11385_ = \bapg_rd.w_ptr_r [1] ? _11384_ : _11383_;
  assign _11386_ = \bapg_rd.w_ptr_r [2] ? _11385_ : _11382_;
  assign _11387_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [10] : \MSYNC_1r1w.synth.nz.mem[88] [10];
  assign _11388_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [10] : \MSYNC_1r1w.synth.nz.mem[90] [10];
  assign _11389_ = \bapg_rd.w_ptr_r [1] ? _11388_ : _11387_;
  assign _11390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [10] : \MSYNC_1r1w.synth.nz.mem[92] [10];
  assign _11391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [10] : \MSYNC_1r1w.synth.nz.mem[94] [10];
  assign _11392_ = \bapg_rd.w_ptr_r [1] ? _11391_ : _11390_;
  assign _11393_ = \bapg_rd.w_ptr_r [2] ? _11392_ : _11389_;
  assign _11394_ = \bapg_rd.w_ptr_r [3] ? _11393_ : _11386_;
  assign _11395_ = \bapg_rd.w_ptr_r [4] ? _11394_ : _11379_;
  assign _11396_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [10] : \MSYNC_1r1w.synth.nz.mem[96] [10];
  assign _11397_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [10] : \MSYNC_1r1w.synth.nz.mem[98] [10];
  assign _11398_ = \bapg_rd.w_ptr_r [1] ? _11397_ : _11396_;
  assign _11399_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [10] : \MSYNC_1r1w.synth.nz.mem[100] [10];
  assign _11400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [10] : \MSYNC_1r1w.synth.nz.mem[102] [10];
  assign _11401_ = \bapg_rd.w_ptr_r [1] ? _11400_ : _11399_;
  assign _11402_ = \bapg_rd.w_ptr_r [2] ? _11401_ : _11398_;
  assign _11403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [10] : \MSYNC_1r1w.synth.nz.mem[104] [10];
  assign _11404_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [10] : \MSYNC_1r1w.synth.nz.mem[106] [10];
  assign _11405_ = \bapg_rd.w_ptr_r [1] ? _11404_ : _11403_;
  assign _11406_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [10] : \MSYNC_1r1w.synth.nz.mem[108] [10];
  assign _11407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [10] : \MSYNC_1r1w.synth.nz.mem[110] [10];
  assign _11408_ = \bapg_rd.w_ptr_r [1] ? _11407_ : _11406_;
  assign _11409_ = \bapg_rd.w_ptr_r [2] ? _11408_ : _11405_;
  assign _11410_ = \bapg_rd.w_ptr_r [3] ? _11409_ : _11402_;
  assign _11411_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [10] : \MSYNC_1r1w.synth.nz.mem[112] [10];
  assign _11412_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [10] : \MSYNC_1r1w.synth.nz.mem[114] [10];
  assign _11413_ = \bapg_rd.w_ptr_r [1] ? _11412_ : _11411_;
  assign _11414_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [10] : \MSYNC_1r1w.synth.nz.mem[116] [10];
  assign _11415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [10] : \MSYNC_1r1w.synth.nz.mem[118] [10];
  assign _11416_ = \bapg_rd.w_ptr_r [1] ? _11415_ : _11414_;
  assign _11417_ = \bapg_rd.w_ptr_r [2] ? _11416_ : _11413_;
  assign _11418_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [10] : \MSYNC_1r1w.synth.nz.mem[120] [10];
  assign _11419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [10] : \MSYNC_1r1w.synth.nz.mem[122] [10];
  assign _11420_ = \bapg_rd.w_ptr_r [1] ? _11419_ : _11418_;
  assign _11421_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [10] : \MSYNC_1r1w.synth.nz.mem[124] [10];
  assign _11422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [10] : \MSYNC_1r1w.synth.nz.mem[126] [10];
  assign _11423_ = \bapg_rd.w_ptr_r [1] ? _11422_ : _11421_;
  assign _11424_ = \bapg_rd.w_ptr_r [2] ? _11423_ : _11420_;
  assign _11425_ = \bapg_rd.w_ptr_r [3] ? _11424_ : _11417_;
  assign _11426_ = \bapg_rd.w_ptr_r [4] ? _11425_ : _11410_;
  assign _11427_ = \bapg_rd.w_ptr_r [5] ? _11426_ : _11395_;
  assign _11428_ = \bapg_rd.w_ptr_r [6] ? _11427_ : _11364_;
  assign _11429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [10] : \MSYNC_1r1w.synth.nz.mem[128] [10];
  assign _11430_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [10] : \MSYNC_1r1w.synth.nz.mem[130] [10];
  assign _11431_ = \bapg_rd.w_ptr_r [1] ? _11430_ : _11429_;
  assign _11432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [10] : \MSYNC_1r1w.synth.nz.mem[132] [10];
  assign _11433_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [10] : \MSYNC_1r1w.synth.nz.mem[134] [10];
  assign _11434_ = \bapg_rd.w_ptr_r [1] ? _11433_ : _11432_;
  assign _11435_ = \bapg_rd.w_ptr_r [2] ? _11434_ : _11431_;
  assign _11436_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [10] : \MSYNC_1r1w.synth.nz.mem[136] [10];
  assign _11437_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [10] : \MSYNC_1r1w.synth.nz.mem[138] [10];
  assign _11438_ = \bapg_rd.w_ptr_r [1] ? _11437_ : _11436_;
  assign _11439_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [10] : \MSYNC_1r1w.synth.nz.mem[140] [10];
  assign _11440_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [10] : \MSYNC_1r1w.synth.nz.mem[142] [10];
  assign _11441_ = \bapg_rd.w_ptr_r [1] ? _11440_ : _11439_;
  assign _11442_ = \bapg_rd.w_ptr_r [2] ? _11441_ : _11438_;
  assign _11443_ = \bapg_rd.w_ptr_r [3] ? _11442_ : _11435_;
  assign _11444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [10] : \MSYNC_1r1w.synth.nz.mem[144] [10];
  assign _11445_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [10] : \MSYNC_1r1w.synth.nz.mem[146] [10];
  assign _11446_ = \bapg_rd.w_ptr_r [1] ? _11445_ : _11444_;
  assign _11447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [10] : \MSYNC_1r1w.synth.nz.mem[148] [10];
  assign _11448_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [10] : \MSYNC_1r1w.synth.nz.mem[150] [10];
  assign _11449_ = \bapg_rd.w_ptr_r [1] ? _11448_ : _11447_;
  assign _11450_ = \bapg_rd.w_ptr_r [2] ? _11449_ : _11446_;
  assign _11451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [10] : \MSYNC_1r1w.synth.nz.mem[152] [10];
  assign _11452_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [10] : \MSYNC_1r1w.synth.nz.mem[154] [10];
  assign _11453_ = \bapg_rd.w_ptr_r [1] ? _11452_ : _11451_;
  assign _11454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [10] : \MSYNC_1r1w.synth.nz.mem[156] [10];
  assign _11455_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [10] : \MSYNC_1r1w.synth.nz.mem[158] [10];
  assign _11456_ = \bapg_rd.w_ptr_r [1] ? _11455_ : _11454_;
  assign _11457_ = \bapg_rd.w_ptr_r [2] ? _11456_ : _11453_;
  assign _11458_ = \bapg_rd.w_ptr_r [3] ? _11457_ : _11450_;
  assign _11459_ = \bapg_rd.w_ptr_r [4] ? _11458_ : _11443_;
  assign _11460_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [10] : \MSYNC_1r1w.synth.nz.mem[160] [10];
  assign _11461_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [10] : \MSYNC_1r1w.synth.nz.mem[162] [10];
  assign _11462_ = \bapg_rd.w_ptr_r [1] ? _11461_ : _11460_;
  assign _11463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [10] : \MSYNC_1r1w.synth.nz.mem[164] [10];
  assign _11464_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [10] : \MSYNC_1r1w.synth.nz.mem[166] [10];
  assign _11465_ = \bapg_rd.w_ptr_r [1] ? _11464_ : _11463_;
  assign _11466_ = \bapg_rd.w_ptr_r [2] ? _11465_ : _11462_;
  assign _11467_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [10] : \MSYNC_1r1w.synth.nz.mem[168] [10];
  assign _11468_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [10] : \MSYNC_1r1w.synth.nz.mem[170] [10];
  assign _11469_ = \bapg_rd.w_ptr_r [1] ? _11468_ : _11467_;
  assign _11470_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [10] : \MSYNC_1r1w.synth.nz.mem[172] [10];
  assign _11471_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [10] : \MSYNC_1r1w.synth.nz.mem[174] [10];
  assign _11472_ = \bapg_rd.w_ptr_r [1] ? _11471_ : _11470_;
  assign _11473_ = \bapg_rd.w_ptr_r [2] ? _11472_ : _11469_;
  assign _11474_ = \bapg_rd.w_ptr_r [3] ? _11473_ : _11466_;
  assign _11475_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [10] : \MSYNC_1r1w.synth.nz.mem[176] [10];
  assign _11476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [10] : \MSYNC_1r1w.synth.nz.mem[178] [10];
  assign _11477_ = \bapg_rd.w_ptr_r [1] ? _11476_ : _11475_;
  assign _11478_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [10] : \MSYNC_1r1w.synth.nz.mem[180] [10];
  assign _11479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [10] : \MSYNC_1r1w.synth.nz.mem[182] [10];
  assign _11480_ = \bapg_rd.w_ptr_r [1] ? _11479_ : _11478_;
  assign _11481_ = \bapg_rd.w_ptr_r [2] ? _11480_ : _11477_;
  assign _11482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [10] : \MSYNC_1r1w.synth.nz.mem[184] [10];
  assign _11483_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [10] : \MSYNC_1r1w.synth.nz.mem[186] [10];
  assign _11484_ = \bapg_rd.w_ptr_r [1] ? _11483_ : _11482_;
  assign _11485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [10] : \MSYNC_1r1w.synth.nz.mem[188] [10];
  assign _11486_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [10] : \MSYNC_1r1w.synth.nz.mem[190] [10];
  assign _11487_ = \bapg_rd.w_ptr_r [1] ? _11486_ : _11485_;
  assign _11488_ = \bapg_rd.w_ptr_r [2] ? _11487_ : _11484_;
  assign _11489_ = \bapg_rd.w_ptr_r [3] ? _11488_ : _11481_;
  assign _11490_ = \bapg_rd.w_ptr_r [4] ? _11489_ : _11474_;
  assign _11491_ = \bapg_rd.w_ptr_r [5] ? _11490_ : _11459_;
  assign _11492_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [10] : \MSYNC_1r1w.synth.nz.mem[192] [10];
  assign _11493_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [10] : \MSYNC_1r1w.synth.nz.mem[194] [10];
  assign _11494_ = \bapg_rd.w_ptr_r [1] ? _11493_ : _11492_;
  assign _11495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [10] : \MSYNC_1r1w.synth.nz.mem[196] [10];
  assign _11496_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [10] : \MSYNC_1r1w.synth.nz.mem[198] [10];
  assign _11497_ = \bapg_rd.w_ptr_r [1] ? _11496_ : _11495_;
  assign _11498_ = \bapg_rd.w_ptr_r [2] ? _11497_ : _11494_;
  assign _11499_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [10] : \MSYNC_1r1w.synth.nz.mem[200] [10];
  assign _11500_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [10] : \MSYNC_1r1w.synth.nz.mem[202] [10];
  assign _11501_ = \bapg_rd.w_ptr_r [1] ? _11500_ : _11499_;
  assign _11502_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [10] : \MSYNC_1r1w.synth.nz.mem[204] [10];
  assign _11503_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [10] : \MSYNC_1r1w.synth.nz.mem[206] [10];
  assign _11504_ = \bapg_rd.w_ptr_r [1] ? _11503_ : _11502_;
  assign _11505_ = \bapg_rd.w_ptr_r [2] ? _11504_ : _11501_;
  assign _11506_ = \bapg_rd.w_ptr_r [3] ? _11505_ : _11498_;
  assign _11507_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [10] : \MSYNC_1r1w.synth.nz.mem[208] [10];
  assign _11508_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [10] : \MSYNC_1r1w.synth.nz.mem[210] [10];
  assign _11509_ = \bapg_rd.w_ptr_r [1] ? _11508_ : _11507_;
  assign _11510_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [10] : \MSYNC_1r1w.synth.nz.mem[212] [10];
  assign _11511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [10] : \MSYNC_1r1w.synth.nz.mem[214] [10];
  assign _11512_ = \bapg_rd.w_ptr_r [1] ? _11511_ : _11510_;
  assign _11513_ = \bapg_rd.w_ptr_r [2] ? _11512_ : _11509_;
  assign _11514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [10] : \MSYNC_1r1w.synth.nz.mem[216] [10];
  assign _11515_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [10] : \MSYNC_1r1w.synth.nz.mem[218] [10];
  assign _11516_ = \bapg_rd.w_ptr_r [1] ? _11515_ : _11514_;
  assign _11517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [10] : \MSYNC_1r1w.synth.nz.mem[220] [10];
  assign _11518_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [10] : \MSYNC_1r1w.synth.nz.mem[222] [10];
  assign _11519_ = \bapg_rd.w_ptr_r [1] ? _11518_ : _11517_;
  assign _11520_ = \bapg_rd.w_ptr_r [2] ? _11519_ : _11516_;
  assign _11521_ = \bapg_rd.w_ptr_r [3] ? _11520_ : _11513_;
  assign _11522_ = \bapg_rd.w_ptr_r [4] ? _11521_ : _11506_;
  assign _11523_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [10] : \MSYNC_1r1w.synth.nz.mem[224] [10];
  assign _11524_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [10] : \MSYNC_1r1w.synth.nz.mem[226] [10];
  assign _11525_ = \bapg_rd.w_ptr_r [1] ? _11524_ : _11523_;
  assign _11526_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [10] : \MSYNC_1r1w.synth.nz.mem[228] [10];
  assign _11527_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [10] : \MSYNC_1r1w.synth.nz.mem[230] [10];
  assign _11528_ = \bapg_rd.w_ptr_r [1] ? _11527_ : _11526_;
  assign _11529_ = \bapg_rd.w_ptr_r [2] ? _11528_ : _11525_;
  assign _11530_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [10] : \MSYNC_1r1w.synth.nz.mem[232] [10];
  assign _11531_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [10] : \MSYNC_1r1w.synth.nz.mem[234] [10];
  assign _11532_ = \bapg_rd.w_ptr_r [1] ? _11531_ : _11530_;
  assign _11533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [10] : \MSYNC_1r1w.synth.nz.mem[236] [10];
  assign _11534_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [10] : \MSYNC_1r1w.synth.nz.mem[238] [10];
  assign _11535_ = \bapg_rd.w_ptr_r [1] ? _11534_ : _11533_;
  assign _11536_ = \bapg_rd.w_ptr_r [2] ? _11535_ : _11532_;
  assign _11537_ = \bapg_rd.w_ptr_r [3] ? _11536_ : _11529_;
  assign _11538_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [10] : \MSYNC_1r1w.synth.nz.mem[240] [10];
  assign _11539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [10] : \MSYNC_1r1w.synth.nz.mem[242] [10];
  assign _11540_ = \bapg_rd.w_ptr_r [1] ? _11539_ : _11538_;
  assign _11541_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [10] : \MSYNC_1r1w.synth.nz.mem[244] [10];
  assign _11542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [10] : \MSYNC_1r1w.synth.nz.mem[246] [10];
  assign _11543_ = \bapg_rd.w_ptr_r [1] ? _11542_ : _11541_;
  assign _11544_ = \bapg_rd.w_ptr_r [2] ? _11543_ : _11540_;
  assign _11545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [10] : \MSYNC_1r1w.synth.nz.mem[248] [10];
  assign _11546_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [10] : \MSYNC_1r1w.synth.nz.mem[250] [10];
  assign _11547_ = \bapg_rd.w_ptr_r [1] ? _11546_ : _11545_;
  assign _11548_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [10] : \MSYNC_1r1w.synth.nz.mem[252] [10];
  assign _11549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [10] : \MSYNC_1r1w.synth.nz.mem[254] [10];
  assign _11550_ = \bapg_rd.w_ptr_r [1] ? _11549_ : _11548_;
  assign _11551_ = \bapg_rd.w_ptr_r [2] ? _11550_ : _11547_;
  assign _11552_ = \bapg_rd.w_ptr_r [3] ? _11551_ : _11544_;
  assign _11553_ = \bapg_rd.w_ptr_r [4] ? _11552_ : _11537_;
  assign _11554_ = \bapg_rd.w_ptr_r [5] ? _11553_ : _11522_;
  assign _11555_ = \bapg_rd.w_ptr_r [6] ? _11554_ : _11491_;
  assign _11556_ = \bapg_rd.w_ptr_r [7] ? _11555_ : _11428_;
  assign _11557_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [10] : \MSYNC_1r1w.synth.nz.mem[256] [10];
  assign _11558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [10] : \MSYNC_1r1w.synth.nz.mem[258] [10];
  assign _11559_ = \bapg_rd.w_ptr_r [1] ? _11558_ : _11557_;
  assign _11560_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [10] : \MSYNC_1r1w.synth.nz.mem[260] [10];
  assign _11561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [10] : \MSYNC_1r1w.synth.nz.mem[262] [10];
  assign _11562_ = \bapg_rd.w_ptr_r [1] ? _11561_ : _11560_;
  assign _11563_ = \bapg_rd.w_ptr_r [2] ? _11562_ : _11559_;
  assign _11564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [10] : \MSYNC_1r1w.synth.nz.mem[264] [10];
  assign _11565_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [10] : \MSYNC_1r1w.synth.nz.mem[266] [10];
  assign _11566_ = \bapg_rd.w_ptr_r [1] ? _11565_ : _11564_;
  assign _11567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [10] : \MSYNC_1r1w.synth.nz.mem[268] [10];
  assign _11568_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [10] : \MSYNC_1r1w.synth.nz.mem[270] [10];
  assign _11569_ = \bapg_rd.w_ptr_r [1] ? _11568_ : _11567_;
  assign _11570_ = \bapg_rd.w_ptr_r [2] ? _11569_ : _11566_;
  assign _11571_ = \bapg_rd.w_ptr_r [3] ? _11570_ : _11563_;
  assign _11572_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [10] : \MSYNC_1r1w.synth.nz.mem[272] [10];
  assign _11573_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [10] : \MSYNC_1r1w.synth.nz.mem[274] [10];
  assign _11574_ = \bapg_rd.w_ptr_r [1] ? _11573_ : _11572_;
  assign _11575_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [10] : \MSYNC_1r1w.synth.nz.mem[276] [10];
  assign _11576_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [10] : \MSYNC_1r1w.synth.nz.mem[278] [10];
  assign _11577_ = \bapg_rd.w_ptr_r [1] ? _11576_ : _11575_;
  assign _11578_ = \bapg_rd.w_ptr_r [2] ? _11577_ : _11574_;
  assign _11579_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [10] : \MSYNC_1r1w.synth.nz.mem[280] [10];
  assign _11580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [10] : \MSYNC_1r1w.synth.nz.mem[282] [10];
  assign _11581_ = \bapg_rd.w_ptr_r [1] ? _11580_ : _11579_;
  assign _11582_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [10] : \MSYNC_1r1w.synth.nz.mem[284] [10];
  assign _11583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [10] : \MSYNC_1r1w.synth.nz.mem[286] [10];
  assign _11584_ = \bapg_rd.w_ptr_r [1] ? _11583_ : _11582_;
  assign _11585_ = \bapg_rd.w_ptr_r [2] ? _11584_ : _11581_;
  assign _11586_ = \bapg_rd.w_ptr_r [3] ? _11585_ : _11578_;
  assign _11587_ = \bapg_rd.w_ptr_r [4] ? _11586_ : _11571_;
  assign _11588_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [10] : \MSYNC_1r1w.synth.nz.mem[288] [10];
  assign _11589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [10] : \MSYNC_1r1w.synth.nz.mem[290] [10];
  assign _11590_ = \bapg_rd.w_ptr_r [1] ? _11589_ : _11588_;
  assign _11591_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [10] : \MSYNC_1r1w.synth.nz.mem[292] [10];
  assign _11592_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [10] : \MSYNC_1r1w.synth.nz.mem[294] [10];
  assign _11593_ = \bapg_rd.w_ptr_r [1] ? _11592_ : _11591_;
  assign _11594_ = \bapg_rd.w_ptr_r [2] ? _11593_ : _11590_;
  assign _11595_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [10] : \MSYNC_1r1w.synth.nz.mem[296] [10];
  assign _11596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [10] : \MSYNC_1r1w.synth.nz.mem[298] [10];
  assign _11597_ = \bapg_rd.w_ptr_r [1] ? _11596_ : _11595_;
  assign _11598_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [10] : \MSYNC_1r1w.synth.nz.mem[300] [10];
  assign _11599_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [10] : \MSYNC_1r1w.synth.nz.mem[302] [10];
  assign _11600_ = \bapg_rd.w_ptr_r [1] ? _11599_ : _11598_;
  assign _11601_ = \bapg_rd.w_ptr_r [2] ? _11600_ : _11597_;
  assign _11602_ = \bapg_rd.w_ptr_r [3] ? _11601_ : _11594_;
  assign _11603_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [10] : \MSYNC_1r1w.synth.nz.mem[304] [10];
  assign _11604_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [10] : \MSYNC_1r1w.synth.nz.mem[306] [10];
  assign _11605_ = \bapg_rd.w_ptr_r [1] ? _11604_ : _11603_;
  assign _11606_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [10] : \MSYNC_1r1w.synth.nz.mem[308] [10];
  assign _11607_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [10] : \MSYNC_1r1w.synth.nz.mem[310] [10];
  assign _11608_ = \bapg_rd.w_ptr_r [1] ? _11607_ : _11606_;
  assign _11609_ = \bapg_rd.w_ptr_r [2] ? _11608_ : _11605_;
  assign _11610_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [10] : \MSYNC_1r1w.synth.nz.mem[312] [10];
  assign _11611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [10] : \MSYNC_1r1w.synth.nz.mem[314] [10];
  assign _11612_ = \bapg_rd.w_ptr_r [1] ? _11611_ : _11610_;
  assign _11613_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [10] : \MSYNC_1r1w.synth.nz.mem[316] [10];
  assign _11614_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [10] : \MSYNC_1r1w.synth.nz.mem[318] [10];
  assign _11615_ = \bapg_rd.w_ptr_r [1] ? _11614_ : _11613_;
  assign _11616_ = \bapg_rd.w_ptr_r [2] ? _11615_ : _11612_;
  assign _11617_ = \bapg_rd.w_ptr_r [3] ? _11616_ : _11609_;
  assign _11618_ = \bapg_rd.w_ptr_r [4] ? _11617_ : _11602_;
  assign _11619_ = \bapg_rd.w_ptr_r [5] ? _11618_ : _11587_;
  assign _11620_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [10] : \MSYNC_1r1w.synth.nz.mem[320] [10];
  assign _11621_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [10] : \MSYNC_1r1w.synth.nz.mem[322] [10];
  assign _11622_ = \bapg_rd.w_ptr_r [1] ? _11621_ : _11620_;
  assign _11623_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [10] : \MSYNC_1r1w.synth.nz.mem[324] [10];
  assign _11624_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [10] : \MSYNC_1r1w.synth.nz.mem[326] [10];
  assign _11625_ = \bapg_rd.w_ptr_r [1] ? _11624_ : _11623_;
  assign _11626_ = \bapg_rd.w_ptr_r [2] ? _11625_ : _11622_;
  assign _11627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [10] : \MSYNC_1r1w.synth.nz.mem[328] [10];
  assign _11628_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [10] : \MSYNC_1r1w.synth.nz.mem[330] [10];
  assign _11629_ = \bapg_rd.w_ptr_r [1] ? _11628_ : _11627_;
  assign _11630_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [10] : \MSYNC_1r1w.synth.nz.mem[332] [10];
  assign _11631_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [10] : \MSYNC_1r1w.synth.nz.mem[334] [10];
  assign _11632_ = \bapg_rd.w_ptr_r [1] ? _11631_ : _11630_;
  assign _11633_ = \bapg_rd.w_ptr_r [2] ? _11632_ : _11629_;
  assign _11634_ = \bapg_rd.w_ptr_r [3] ? _11633_ : _11626_;
  assign _11635_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [10] : \MSYNC_1r1w.synth.nz.mem[336] [10];
  assign _11636_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [10] : \MSYNC_1r1w.synth.nz.mem[338] [10];
  assign _11637_ = \bapg_rd.w_ptr_r [1] ? _11636_ : _11635_;
  assign _11638_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [10] : \MSYNC_1r1w.synth.nz.mem[340] [10];
  assign _11639_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [10] : \MSYNC_1r1w.synth.nz.mem[342] [10];
  assign _11640_ = \bapg_rd.w_ptr_r [1] ? _11639_ : _11638_;
  assign _11641_ = \bapg_rd.w_ptr_r [2] ? _11640_ : _11637_;
  assign _11642_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [10] : \MSYNC_1r1w.synth.nz.mem[344] [10];
  assign _11643_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [10] : \MSYNC_1r1w.synth.nz.mem[346] [10];
  assign _11644_ = \bapg_rd.w_ptr_r [1] ? _11643_ : _11642_;
  assign _11645_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [10] : \MSYNC_1r1w.synth.nz.mem[348] [10];
  assign _11646_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [10] : \MSYNC_1r1w.synth.nz.mem[350] [10];
  assign _11647_ = \bapg_rd.w_ptr_r [1] ? _11646_ : _11645_;
  assign _11648_ = \bapg_rd.w_ptr_r [2] ? _11647_ : _11644_;
  assign _11649_ = \bapg_rd.w_ptr_r [3] ? _11648_ : _11641_;
  assign _11650_ = \bapg_rd.w_ptr_r [4] ? _11649_ : _11634_;
  assign _11651_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [10] : \MSYNC_1r1w.synth.nz.mem[352] [10];
  assign _11652_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [10] : \MSYNC_1r1w.synth.nz.mem[354] [10];
  assign _11653_ = \bapg_rd.w_ptr_r [1] ? _11652_ : _11651_;
  assign _11654_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [10] : \MSYNC_1r1w.synth.nz.mem[356] [10];
  assign _11655_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [10] : \MSYNC_1r1w.synth.nz.mem[358] [10];
  assign _11656_ = \bapg_rd.w_ptr_r [1] ? _11655_ : _11654_;
  assign _11657_ = \bapg_rd.w_ptr_r [2] ? _11656_ : _11653_;
  assign _11658_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [10] : \MSYNC_1r1w.synth.nz.mem[360] [10];
  assign _11659_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [10] : \MSYNC_1r1w.synth.nz.mem[362] [10];
  assign _11660_ = \bapg_rd.w_ptr_r [1] ? _11659_ : _11658_;
  assign _11661_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [10] : \MSYNC_1r1w.synth.nz.mem[364] [10];
  assign _11662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [10] : \MSYNC_1r1w.synth.nz.mem[366] [10];
  assign _11663_ = \bapg_rd.w_ptr_r [1] ? _11662_ : _11661_;
  assign _11664_ = \bapg_rd.w_ptr_r [2] ? _11663_ : _11660_;
  assign _11665_ = \bapg_rd.w_ptr_r [3] ? _11664_ : _11657_;
  assign _11666_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [10] : \MSYNC_1r1w.synth.nz.mem[368] [10];
  assign _11667_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [10] : \MSYNC_1r1w.synth.nz.mem[370] [10];
  assign _11668_ = \bapg_rd.w_ptr_r [1] ? _11667_ : _11666_;
  assign _11669_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [10] : \MSYNC_1r1w.synth.nz.mem[372] [10];
  assign _11670_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [10] : \MSYNC_1r1w.synth.nz.mem[374] [10];
  assign _11671_ = \bapg_rd.w_ptr_r [1] ? _11670_ : _11669_;
  assign _11672_ = \bapg_rd.w_ptr_r [2] ? _11671_ : _11668_;
  assign _11673_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [10] : \MSYNC_1r1w.synth.nz.mem[376] [10];
  assign _11674_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [10] : \MSYNC_1r1w.synth.nz.mem[378] [10];
  assign _11675_ = \bapg_rd.w_ptr_r [1] ? _11674_ : _11673_;
  assign _11676_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [10] : \MSYNC_1r1w.synth.nz.mem[380] [10];
  assign _11677_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [10] : \MSYNC_1r1w.synth.nz.mem[382] [10];
  assign _11678_ = \bapg_rd.w_ptr_r [1] ? _11677_ : _11676_;
  assign _11679_ = \bapg_rd.w_ptr_r [2] ? _11678_ : _11675_;
  assign _11680_ = \bapg_rd.w_ptr_r [3] ? _11679_ : _11672_;
  assign _11681_ = \bapg_rd.w_ptr_r [4] ? _11680_ : _11665_;
  assign _11682_ = \bapg_rd.w_ptr_r [5] ? _11681_ : _11650_;
  assign _11683_ = \bapg_rd.w_ptr_r [6] ? _11682_ : _11619_;
  assign _11684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [10] : \MSYNC_1r1w.synth.nz.mem[384] [10];
  assign _11685_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [10] : \MSYNC_1r1w.synth.nz.mem[386] [10];
  assign _11686_ = \bapg_rd.w_ptr_r [1] ? _11685_ : _11684_;
  assign _11687_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [10] : \MSYNC_1r1w.synth.nz.mem[388] [10];
  assign _11688_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [10] : \MSYNC_1r1w.synth.nz.mem[390] [10];
  assign _11689_ = \bapg_rd.w_ptr_r [1] ? _11688_ : _11687_;
  assign _11690_ = \bapg_rd.w_ptr_r [2] ? _11689_ : _11686_;
  assign _11691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [10] : \MSYNC_1r1w.synth.nz.mem[392] [10];
  assign _11692_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [10] : \MSYNC_1r1w.synth.nz.mem[394] [10];
  assign _11693_ = \bapg_rd.w_ptr_r [1] ? _11692_ : _11691_;
  assign _11694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [10] : \MSYNC_1r1w.synth.nz.mem[396] [10];
  assign _11695_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [10] : \MSYNC_1r1w.synth.nz.mem[398] [10];
  assign _11696_ = \bapg_rd.w_ptr_r [1] ? _11695_ : _11694_;
  assign _11697_ = \bapg_rd.w_ptr_r [2] ? _11696_ : _11693_;
  assign _11698_ = \bapg_rd.w_ptr_r [3] ? _11697_ : _11690_;
  assign _11699_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [10] : \MSYNC_1r1w.synth.nz.mem[400] [10];
  assign _11700_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [10] : \MSYNC_1r1w.synth.nz.mem[402] [10];
  assign _11701_ = \bapg_rd.w_ptr_r [1] ? _11700_ : _11699_;
  assign _11702_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [10] : \MSYNC_1r1w.synth.nz.mem[404] [10];
  assign _11703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [10] : \MSYNC_1r1w.synth.nz.mem[406] [10];
  assign _11704_ = \bapg_rd.w_ptr_r [1] ? _11703_ : _11702_;
  assign _11705_ = \bapg_rd.w_ptr_r [2] ? _11704_ : _11701_;
  assign _11706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [10] : \MSYNC_1r1w.synth.nz.mem[408] [10];
  assign _11707_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [10] : \MSYNC_1r1w.synth.nz.mem[410] [10];
  assign _11708_ = \bapg_rd.w_ptr_r [1] ? _11707_ : _11706_;
  assign _11709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [10] : \MSYNC_1r1w.synth.nz.mem[412] [10];
  assign _11710_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [10] : \MSYNC_1r1w.synth.nz.mem[414] [10];
  assign _11711_ = \bapg_rd.w_ptr_r [1] ? _11710_ : _11709_;
  assign _11712_ = \bapg_rd.w_ptr_r [2] ? _11711_ : _11708_;
  assign _11713_ = \bapg_rd.w_ptr_r [3] ? _11712_ : _11705_;
  assign _11714_ = \bapg_rd.w_ptr_r [4] ? _11713_ : _11698_;
  assign _11715_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [10] : \MSYNC_1r1w.synth.nz.mem[416] [10];
  assign _11716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [10] : \MSYNC_1r1w.synth.nz.mem[418] [10];
  assign _11717_ = \bapg_rd.w_ptr_r [1] ? _11716_ : _11715_;
  assign _11718_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [10] : \MSYNC_1r1w.synth.nz.mem[420] [10];
  assign _11719_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [10] : \MSYNC_1r1w.synth.nz.mem[422] [10];
  assign _11720_ = \bapg_rd.w_ptr_r [1] ? _11719_ : _11718_;
  assign _11721_ = \bapg_rd.w_ptr_r [2] ? _11720_ : _11717_;
  assign _11722_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [10] : \MSYNC_1r1w.synth.nz.mem[424] [10];
  assign _11723_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [10] : \MSYNC_1r1w.synth.nz.mem[426] [10];
  assign _11724_ = \bapg_rd.w_ptr_r [1] ? _11723_ : _11722_;
  assign _11725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [10] : \MSYNC_1r1w.synth.nz.mem[428] [10];
  assign _11726_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [10] : \MSYNC_1r1w.synth.nz.mem[430] [10];
  assign _11727_ = \bapg_rd.w_ptr_r [1] ? _11726_ : _11725_;
  assign _11728_ = \bapg_rd.w_ptr_r [2] ? _11727_ : _11724_;
  assign _11729_ = \bapg_rd.w_ptr_r [3] ? _11728_ : _11721_;
  assign _11730_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [10] : \MSYNC_1r1w.synth.nz.mem[432] [10];
  assign _11731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [10] : \MSYNC_1r1w.synth.nz.mem[434] [10];
  assign _11732_ = \bapg_rd.w_ptr_r [1] ? _11731_ : _11730_;
  assign _11733_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [10] : \MSYNC_1r1w.synth.nz.mem[436] [10];
  assign _11734_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [10] : \MSYNC_1r1w.synth.nz.mem[438] [10];
  assign _11735_ = \bapg_rd.w_ptr_r [1] ? _11734_ : _11733_;
  assign _11736_ = \bapg_rd.w_ptr_r [2] ? _11735_ : _11732_;
  assign _11737_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [10] : \MSYNC_1r1w.synth.nz.mem[440] [10];
  assign _11738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [10] : \MSYNC_1r1w.synth.nz.mem[442] [10];
  assign _11739_ = \bapg_rd.w_ptr_r [1] ? _11738_ : _11737_;
  assign _11740_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [10] : \MSYNC_1r1w.synth.nz.mem[444] [10];
  assign _11741_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [10] : \MSYNC_1r1w.synth.nz.mem[446] [10];
  assign _11742_ = \bapg_rd.w_ptr_r [1] ? _11741_ : _11740_;
  assign _11743_ = \bapg_rd.w_ptr_r [2] ? _11742_ : _11739_;
  assign _11744_ = \bapg_rd.w_ptr_r [3] ? _11743_ : _11736_;
  assign _11745_ = \bapg_rd.w_ptr_r [4] ? _11744_ : _11729_;
  assign _11746_ = \bapg_rd.w_ptr_r [5] ? _11745_ : _11714_;
  assign _11747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [10] : \MSYNC_1r1w.synth.nz.mem[448] [10];
  assign _11748_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [10] : \MSYNC_1r1w.synth.nz.mem[450] [10];
  assign _11749_ = \bapg_rd.w_ptr_r [1] ? _11748_ : _11747_;
  assign _11750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [10] : \MSYNC_1r1w.synth.nz.mem[452] [10];
  assign _11751_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [10] : \MSYNC_1r1w.synth.nz.mem[454] [10];
  assign _11752_ = \bapg_rd.w_ptr_r [1] ? _11751_ : _11750_;
  assign _11753_ = \bapg_rd.w_ptr_r [2] ? _11752_ : _11749_;
  assign _11754_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [10] : \MSYNC_1r1w.synth.nz.mem[456] [10];
  assign _11755_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [10] : \MSYNC_1r1w.synth.nz.mem[458] [10];
  assign _11756_ = \bapg_rd.w_ptr_r [1] ? _11755_ : _11754_;
  assign _11757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [10] : \MSYNC_1r1w.synth.nz.mem[460] [10];
  assign _11758_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [10] : \MSYNC_1r1w.synth.nz.mem[462] [10];
  assign _11759_ = \bapg_rd.w_ptr_r [1] ? _11758_ : _11757_;
  assign _11760_ = \bapg_rd.w_ptr_r [2] ? _11759_ : _11756_;
  assign _11761_ = \bapg_rd.w_ptr_r [3] ? _11760_ : _11753_;
  assign _11762_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [10] : \MSYNC_1r1w.synth.nz.mem[464] [10];
  assign _11763_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [10] : \MSYNC_1r1w.synth.nz.mem[466] [10];
  assign _11764_ = \bapg_rd.w_ptr_r [1] ? _11763_ : _11762_;
  assign _11765_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [10] : \MSYNC_1r1w.synth.nz.mem[468] [10];
  assign _11766_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [10] : \MSYNC_1r1w.synth.nz.mem[470] [10];
  assign _11767_ = \bapg_rd.w_ptr_r [1] ? _11766_ : _11765_;
  assign _11768_ = \bapg_rd.w_ptr_r [2] ? _11767_ : _11764_;
  assign _11769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [10] : \MSYNC_1r1w.synth.nz.mem[472] [10];
  assign _11770_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [10] : \MSYNC_1r1w.synth.nz.mem[474] [10];
  assign _11771_ = \bapg_rd.w_ptr_r [1] ? _11770_ : _11769_;
  assign _11772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [10] : \MSYNC_1r1w.synth.nz.mem[476] [10];
  assign _11773_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [10] : \MSYNC_1r1w.synth.nz.mem[478] [10];
  assign _11774_ = \bapg_rd.w_ptr_r [1] ? _11773_ : _11772_;
  assign _11775_ = \bapg_rd.w_ptr_r [2] ? _11774_ : _11771_;
  assign _11776_ = \bapg_rd.w_ptr_r [3] ? _11775_ : _11768_;
  assign _11777_ = \bapg_rd.w_ptr_r [4] ? _11776_ : _11761_;
  assign _11778_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [10] : \MSYNC_1r1w.synth.nz.mem[480] [10];
  assign _11779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [10] : \MSYNC_1r1w.synth.nz.mem[482] [10];
  assign _11780_ = \bapg_rd.w_ptr_r [1] ? _11779_ : _11778_;
  assign _11781_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [10] : \MSYNC_1r1w.synth.nz.mem[484] [10];
  assign _11782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [10] : \MSYNC_1r1w.synth.nz.mem[486] [10];
  assign _11783_ = \bapg_rd.w_ptr_r [1] ? _11782_ : _11781_;
  assign _11784_ = \bapg_rd.w_ptr_r [2] ? _11783_ : _11780_;
  assign _11785_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [10] : \MSYNC_1r1w.synth.nz.mem[488] [10];
  assign _11786_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [10] : \MSYNC_1r1w.synth.nz.mem[490] [10];
  assign _11787_ = \bapg_rd.w_ptr_r [1] ? _11786_ : _11785_;
  assign _11788_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [10] : \MSYNC_1r1w.synth.nz.mem[492] [10];
  assign _11789_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [10] : \MSYNC_1r1w.synth.nz.mem[494] [10];
  assign _11790_ = \bapg_rd.w_ptr_r [1] ? _11789_ : _11788_;
  assign _11791_ = \bapg_rd.w_ptr_r [2] ? _11790_ : _11787_;
  assign _11792_ = \bapg_rd.w_ptr_r [3] ? _11791_ : _11784_;
  assign _11793_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [10] : \MSYNC_1r1w.synth.nz.mem[496] [10];
  assign _11794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [10] : \MSYNC_1r1w.synth.nz.mem[498] [10];
  assign _11795_ = \bapg_rd.w_ptr_r [1] ? _11794_ : _11793_;
  assign _11796_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [10] : \MSYNC_1r1w.synth.nz.mem[500] [10];
  assign _11797_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [10] : \MSYNC_1r1w.synth.nz.mem[502] [10];
  assign _11798_ = \bapg_rd.w_ptr_r [1] ? _11797_ : _11796_;
  assign _11799_ = \bapg_rd.w_ptr_r [2] ? _11798_ : _11795_;
  assign _11800_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [10] : \MSYNC_1r1w.synth.nz.mem[504] [10];
  assign _11801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [10] : \MSYNC_1r1w.synth.nz.mem[506] [10];
  assign _11802_ = \bapg_rd.w_ptr_r [1] ? _11801_ : _11800_;
  assign _11803_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [10] : \MSYNC_1r1w.synth.nz.mem[508] [10];
  assign _11804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [10] : \MSYNC_1r1w.synth.nz.mem[510] [10];
  assign _11805_ = \bapg_rd.w_ptr_r [1] ? _11804_ : _11803_;
  assign _11806_ = \bapg_rd.w_ptr_r [2] ? _11805_ : _11802_;
  assign _11807_ = \bapg_rd.w_ptr_r [3] ? _11806_ : _11799_;
  assign _11808_ = \bapg_rd.w_ptr_r [4] ? _11807_ : _11792_;
  assign _11809_ = \bapg_rd.w_ptr_r [5] ? _11808_ : _11777_;
  assign _11810_ = \bapg_rd.w_ptr_r [6] ? _11809_ : _11746_;
  assign _11811_ = \bapg_rd.w_ptr_r [7] ? _11810_ : _11683_;
  assign _11812_ = \bapg_rd.w_ptr_r [8] ? _11811_ : _11556_;
  assign _11813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [10] : \MSYNC_1r1w.synth.nz.mem[512] [10];
  assign _11814_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [10] : \MSYNC_1r1w.synth.nz.mem[514] [10];
  assign _11815_ = \bapg_rd.w_ptr_r [1] ? _11814_ : _11813_;
  assign _11816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [10] : \MSYNC_1r1w.synth.nz.mem[516] [10];
  assign _11817_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [10] : \MSYNC_1r1w.synth.nz.mem[518] [10];
  assign _11818_ = \bapg_rd.w_ptr_r [1] ? _11817_ : _11816_;
  assign _11819_ = \bapg_rd.w_ptr_r [2] ? _11818_ : _11815_;
  assign _11820_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [10] : \MSYNC_1r1w.synth.nz.mem[520] [10];
  assign _11821_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [10] : \MSYNC_1r1w.synth.nz.mem[522] [10];
  assign _11822_ = \bapg_rd.w_ptr_r [1] ? _11821_ : _11820_;
  assign _11823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [10] : \MSYNC_1r1w.synth.nz.mem[524] [10];
  assign _11824_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [10] : \MSYNC_1r1w.synth.nz.mem[526] [10];
  assign _11825_ = \bapg_rd.w_ptr_r [1] ? _11824_ : _11823_;
  assign _11826_ = \bapg_rd.w_ptr_r [2] ? _11825_ : _11822_;
  assign _11827_ = \bapg_rd.w_ptr_r [3] ? _11826_ : _11819_;
  assign _11828_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [10] : \MSYNC_1r1w.synth.nz.mem[528] [10];
  assign _11829_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [10] : \MSYNC_1r1w.synth.nz.mem[530] [10];
  assign _11830_ = \bapg_rd.w_ptr_r [1] ? _11829_ : _11828_;
  assign _11831_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [10] : \MSYNC_1r1w.synth.nz.mem[532] [10];
  assign _11832_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [10] : \MSYNC_1r1w.synth.nz.mem[534] [10];
  assign _11833_ = \bapg_rd.w_ptr_r [1] ? _11832_ : _11831_;
  assign _11834_ = \bapg_rd.w_ptr_r [2] ? _11833_ : _11830_;
  assign _11835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [10] : \MSYNC_1r1w.synth.nz.mem[536] [10];
  assign _11836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [10] : \MSYNC_1r1w.synth.nz.mem[538] [10];
  assign _11837_ = \bapg_rd.w_ptr_r [1] ? _11836_ : _11835_;
  assign _11838_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [10] : \MSYNC_1r1w.synth.nz.mem[540] [10];
  assign _11839_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [10] : \MSYNC_1r1w.synth.nz.mem[542] [10];
  assign _11840_ = \bapg_rd.w_ptr_r [1] ? _11839_ : _11838_;
  assign _11841_ = \bapg_rd.w_ptr_r [2] ? _11840_ : _11837_;
  assign _11842_ = \bapg_rd.w_ptr_r [3] ? _11841_ : _11834_;
  assign _11843_ = \bapg_rd.w_ptr_r [4] ? _11842_ : _11827_;
  assign _11844_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [10] : \MSYNC_1r1w.synth.nz.mem[544] [10];
  assign _11845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [10] : \MSYNC_1r1w.synth.nz.mem[546] [10];
  assign _11846_ = \bapg_rd.w_ptr_r [1] ? _11845_ : _11844_;
  assign _11847_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [10] : \MSYNC_1r1w.synth.nz.mem[548] [10];
  assign _11848_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [10] : \MSYNC_1r1w.synth.nz.mem[550] [10];
  assign _11849_ = \bapg_rd.w_ptr_r [1] ? _11848_ : _11847_;
  assign _11850_ = \bapg_rd.w_ptr_r [2] ? _11849_ : _11846_;
  assign _11851_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [10] : \MSYNC_1r1w.synth.nz.mem[552] [10];
  assign _11852_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [10] : \MSYNC_1r1w.synth.nz.mem[554] [10];
  assign _11853_ = \bapg_rd.w_ptr_r [1] ? _11852_ : _11851_;
  assign _11854_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [10] : \MSYNC_1r1w.synth.nz.mem[556] [10];
  assign _11855_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [10] : \MSYNC_1r1w.synth.nz.mem[558] [10];
  assign _11856_ = \bapg_rd.w_ptr_r [1] ? _11855_ : _11854_;
  assign _11857_ = \bapg_rd.w_ptr_r [2] ? _11856_ : _11853_;
  assign _11858_ = \bapg_rd.w_ptr_r [3] ? _11857_ : _11850_;
  assign _11859_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [10] : \MSYNC_1r1w.synth.nz.mem[560] [10];
  assign _11860_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [10] : \MSYNC_1r1w.synth.nz.mem[562] [10];
  assign _11861_ = \bapg_rd.w_ptr_r [1] ? _11860_ : _11859_;
  assign _11862_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [10] : \MSYNC_1r1w.synth.nz.mem[564] [10];
  assign _11863_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [10] : \MSYNC_1r1w.synth.nz.mem[566] [10];
  assign _11864_ = \bapg_rd.w_ptr_r [1] ? _11863_ : _11862_;
  assign _11865_ = \bapg_rd.w_ptr_r [2] ? _11864_ : _11861_;
  assign _11866_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [10] : \MSYNC_1r1w.synth.nz.mem[568] [10];
  assign _11867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [10] : \MSYNC_1r1w.synth.nz.mem[570] [10];
  assign _11868_ = \bapg_rd.w_ptr_r [1] ? _11867_ : _11866_;
  assign _11869_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [10] : \MSYNC_1r1w.synth.nz.mem[572] [10];
  assign _11870_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [10] : \MSYNC_1r1w.synth.nz.mem[574] [10];
  assign _11871_ = \bapg_rd.w_ptr_r [1] ? _11870_ : _11869_;
  assign _11872_ = \bapg_rd.w_ptr_r [2] ? _11871_ : _11868_;
  assign _11873_ = \bapg_rd.w_ptr_r [3] ? _11872_ : _11865_;
  assign _11874_ = \bapg_rd.w_ptr_r [4] ? _11873_ : _11858_;
  assign _11875_ = \bapg_rd.w_ptr_r [5] ? _11874_ : _11843_;
  assign _11876_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [10] : \MSYNC_1r1w.synth.nz.mem[576] [10];
  assign _11877_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [10] : \MSYNC_1r1w.synth.nz.mem[578] [10];
  assign _11878_ = \bapg_rd.w_ptr_r [1] ? _11877_ : _11876_;
  assign _11879_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [10] : \MSYNC_1r1w.synth.nz.mem[580] [10];
  assign _11880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [10] : \MSYNC_1r1w.synth.nz.mem[582] [10];
  assign _11881_ = \bapg_rd.w_ptr_r [1] ? _11880_ : _11879_;
  assign _11882_ = \bapg_rd.w_ptr_r [2] ? _11881_ : _11878_;
  assign _11883_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [10] : \MSYNC_1r1w.synth.nz.mem[584] [10];
  assign _11884_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [10] : \MSYNC_1r1w.synth.nz.mem[586] [10];
  assign _11885_ = \bapg_rd.w_ptr_r [1] ? _11884_ : _11883_;
  assign _11886_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [10] : \MSYNC_1r1w.synth.nz.mem[588] [10];
  assign _11887_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [10] : \MSYNC_1r1w.synth.nz.mem[590] [10];
  assign _11888_ = \bapg_rd.w_ptr_r [1] ? _11887_ : _11886_;
  assign _11889_ = \bapg_rd.w_ptr_r [2] ? _11888_ : _11885_;
  assign _11890_ = \bapg_rd.w_ptr_r [3] ? _11889_ : _11882_;
  assign _11891_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [10] : \MSYNC_1r1w.synth.nz.mem[592] [10];
  assign _11892_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [10] : \MSYNC_1r1w.synth.nz.mem[594] [10];
  assign _11893_ = \bapg_rd.w_ptr_r [1] ? _11892_ : _11891_;
  assign _11894_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [10] : \MSYNC_1r1w.synth.nz.mem[596] [10];
  assign _11895_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [10] : \MSYNC_1r1w.synth.nz.mem[598] [10];
  assign _11896_ = \bapg_rd.w_ptr_r [1] ? _11895_ : _11894_;
  assign _11897_ = \bapg_rd.w_ptr_r [2] ? _11896_ : _11893_;
  assign _11898_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [10] : \MSYNC_1r1w.synth.nz.mem[600] [10];
  assign _11899_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [10] : \MSYNC_1r1w.synth.nz.mem[602] [10];
  assign _11900_ = \bapg_rd.w_ptr_r [1] ? _11899_ : _11898_;
  assign _11901_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [10] : \MSYNC_1r1w.synth.nz.mem[604] [10];
  assign _11902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [10] : \MSYNC_1r1w.synth.nz.mem[606] [10];
  assign _11903_ = \bapg_rd.w_ptr_r [1] ? _11902_ : _11901_;
  assign _11904_ = \bapg_rd.w_ptr_r [2] ? _11903_ : _11900_;
  assign _11905_ = \bapg_rd.w_ptr_r [3] ? _11904_ : _11897_;
  assign _11906_ = \bapg_rd.w_ptr_r [4] ? _11905_ : _11890_;
  assign _11907_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [10] : \MSYNC_1r1w.synth.nz.mem[608] [10];
  assign _11908_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [10] : \MSYNC_1r1w.synth.nz.mem[610] [10];
  assign _11909_ = \bapg_rd.w_ptr_r [1] ? _11908_ : _11907_;
  assign _11910_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [10] : \MSYNC_1r1w.synth.nz.mem[612] [10];
  assign _11911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [10] : \MSYNC_1r1w.synth.nz.mem[614] [10];
  assign _11912_ = \bapg_rd.w_ptr_r [1] ? _11911_ : _11910_;
  assign _11913_ = \bapg_rd.w_ptr_r [2] ? _11912_ : _11909_;
  assign _11914_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [10] : \MSYNC_1r1w.synth.nz.mem[616] [10];
  assign _11915_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [10] : \MSYNC_1r1w.synth.nz.mem[618] [10];
  assign _11916_ = \bapg_rd.w_ptr_r [1] ? _11915_ : _11914_;
  assign _11917_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [10] : \MSYNC_1r1w.synth.nz.mem[620] [10];
  assign _11918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [10] : \MSYNC_1r1w.synth.nz.mem[622] [10];
  assign _11919_ = \bapg_rd.w_ptr_r [1] ? _11918_ : _11917_;
  assign _11920_ = \bapg_rd.w_ptr_r [2] ? _11919_ : _11916_;
  assign _11921_ = \bapg_rd.w_ptr_r [3] ? _11920_ : _11913_;
  assign _11922_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [10] : \MSYNC_1r1w.synth.nz.mem[624] [10];
  assign _11923_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [10] : \MSYNC_1r1w.synth.nz.mem[626] [10];
  assign _11924_ = \bapg_rd.w_ptr_r [1] ? _11923_ : _11922_;
  assign _11925_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [10] : \MSYNC_1r1w.synth.nz.mem[628] [10];
  assign _11926_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [10] : \MSYNC_1r1w.synth.nz.mem[630] [10];
  assign _11927_ = \bapg_rd.w_ptr_r [1] ? _11926_ : _11925_;
  assign _11928_ = \bapg_rd.w_ptr_r [2] ? _11927_ : _11924_;
  assign _11929_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [10] : \MSYNC_1r1w.synth.nz.mem[632] [10];
  assign _11930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [10] : \MSYNC_1r1w.synth.nz.mem[634] [10];
  assign _11931_ = \bapg_rd.w_ptr_r [1] ? _11930_ : _11929_;
  assign _11932_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [10] : \MSYNC_1r1w.synth.nz.mem[636] [10];
  assign _11933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [10] : \MSYNC_1r1w.synth.nz.mem[638] [10];
  assign _11934_ = \bapg_rd.w_ptr_r [1] ? _11933_ : _11932_;
  assign _11935_ = \bapg_rd.w_ptr_r [2] ? _11934_ : _11931_;
  assign _11936_ = \bapg_rd.w_ptr_r [3] ? _11935_ : _11928_;
  assign _11937_ = \bapg_rd.w_ptr_r [4] ? _11936_ : _11921_;
  assign _11938_ = \bapg_rd.w_ptr_r [5] ? _11937_ : _11906_;
  assign _11939_ = \bapg_rd.w_ptr_r [6] ? _11938_ : _11875_;
  assign _11940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [10] : \MSYNC_1r1w.synth.nz.mem[640] [10];
  assign _11941_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [10] : \MSYNC_1r1w.synth.nz.mem[642] [10];
  assign _11942_ = \bapg_rd.w_ptr_r [1] ? _11941_ : _11940_;
  assign _11943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [10] : \MSYNC_1r1w.synth.nz.mem[644] [10];
  assign _11944_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [10] : \MSYNC_1r1w.synth.nz.mem[646] [10];
  assign _11945_ = \bapg_rd.w_ptr_r [1] ? _11944_ : _11943_;
  assign _11946_ = \bapg_rd.w_ptr_r [2] ? _11945_ : _11942_;
  assign _11947_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [10] : \MSYNC_1r1w.synth.nz.mem[648] [10];
  assign _11948_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [10] : \MSYNC_1r1w.synth.nz.mem[650] [10];
  assign _11949_ = \bapg_rd.w_ptr_r [1] ? _11948_ : _11947_;
  assign _11950_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [10] : \MSYNC_1r1w.synth.nz.mem[652] [10];
  assign _11951_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [10] : \MSYNC_1r1w.synth.nz.mem[654] [10];
  assign _11952_ = \bapg_rd.w_ptr_r [1] ? _11951_ : _11950_;
  assign _11953_ = \bapg_rd.w_ptr_r [2] ? _11952_ : _11949_;
  assign _11954_ = \bapg_rd.w_ptr_r [3] ? _11953_ : _11946_;
  assign _11955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [10] : \MSYNC_1r1w.synth.nz.mem[656] [10];
  assign _11956_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [10] : \MSYNC_1r1w.synth.nz.mem[658] [10];
  assign _11957_ = \bapg_rd.w_ptr_r [1] ? _11956_ : _11955_;
  assign _11958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [10] : \MSYNC_1r1w.synth.nz.mem[660] [10];
  assign _11959_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [10] : \MSYNC_1r1w.synth.nz.mem[662] [10];
  assign _11960_ = \bapg_rd.w_ptr_r [1] ? _11959_ : _11958_;
  assign _11961_ = \bapg_rd.w_ptr_r [2] ? _11960_ : _11957_;
  assign _11962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [10] : \MSYNC_1r1w.synth.nz.mem[664] [10];
  assign _11963_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [10] : \MSYNC_1r1w.synth.nz.mem[666] [10];
  assign _11964_ = \bapg_rd.w_ptr_r [1] ? _11963_ : _11962_;
  assign _11965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [10] : \MSYNC_1r1w.synth.nz.mem[668] [10];
  assign _11966_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [10] : \MSYNC_1r1w.synth.nz.mem[670] [10];
  assign _11967_ = \bapg_rd.w_ptr_r [1] ? _11966_ : _11965_;
  assign _11968_ = \bapg_rd.w_ptr_r [2] ? _11967_ : _11964_;
  assign _11969_ = \bapg_rd.w_ptr_r [3] ? _11968_ : _11961_;
  assign _11970_ = \bapg_rd.w_ptr_r [4] ? _11969_ : _11954_;
  assign _11971_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [10] : \MSYNC_1r1w.synth.nz.mem[672] [10];
  assign _11972_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [10] : \MSYNC_1r1w.synth.nz.mem[674] [10];
  assign _11973_ = \bapg_rd.w_ptr_r [1] ? _11972_ : _11971_;
  assign _11974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [10] : \MSYNC_1r1w.synth.nz.mem[676] [10];
  assign _11975_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [10] : \MSYNC_1r1w.synth.nz.mem[678] [10];
  assign _11976_ = \bapg_rd.w_ptr_r [1] ? _11975_ : _11974_;
  assign _11977_ = \bapg_rd.w_ptr_r [2] ? _11976_ : _11973_;
  assign _11978_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [10] : \MSYNC_1r1w.synth.nz.mem[680] [10];
  assign _11979_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [10] : \MSYNC_1r1w.synth.nz.mem[682] [10];
  assign _11980_ = \bapg_rd.w_ptr_r [1] ? _11979_ : _11978_;
  assign _11981_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [10] : \MSYNC_1r1w.synth.nz.mem[684] [10];
  assign _11982_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [10] : \MSYNC_1r1w.synth.nz.mem[686] [10];
  assign _11983_ = \bapg_rd.w_ptr_r [1] ? _11982_ : _11981_;
  assign _11984_ = \bapg_rd.w_ptr_r [2] ? _11983_ : _11980_;
  assign _11985_ = \bapg_rd.w_ptr_r [3] ? _11984_ : _11977_;
  assign _11986_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [10] : \MSYNC_1r1w.synth.nz.mem[688] [10];
  assign _11987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [10] : \MSYNC_1r1w.synth.nz.mem[690] [10];
  assign _11988_ = \bapg_rd.w_ptr_r [1] ? _11987_ : _11986_;
  assign _11989_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [10] : \MSYNC_1r1w.synth.nz.mem[692] [10];
  assign _11990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [10] : \MSYNC_1r1w.synth.nz.mem[694] [10];
  assign _11991_ = \bapg_rd.w_ptr_r [1] ? _11990_ : _11989_;
  assign _11992_ = \bapg_rd.w_ptr_r [2] ? _11991_ : _11988_;
  assign _11993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [10] : \MSYNC_1r1w.synth.nz.mem[696] [10];
  assign _11994_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [10] : \MSYNC_1r1w.synth.nz.mem[698] [10];
  assign _11995_ = \bapg_rd.w_ptr_r [1] ? _11994_ : _11993_;
  assign _11996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [10] : \MSYNC_1r1w.synth.nz.mem[700] [10];
  assign _11997_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [10] : \MSYNC_1r1w.synth.nz.mem[702] [10];
  assign _11998_ = \bapg_rd.w_ptr_r [1] ? _11997_ : _11996_;
  assign _11999_ = \bapg_rd.w_ptr_r [2] ? _11998_ : _11995_;
  assign _12000_ = \bapg_rd.w_ptr_r [3] ? _11999_ : _11992_;
  assign _12001_ = \bapg_rd.w_ptr_r [4] ? _12000_ : _11985_;
  assign _12002_ = \bapg_rd.w_ptr_r [5] ? _12001_ : _11970_;
  assign _12003_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [10] : \MSYNC_1r1w.synth.nz.mem[704] [10];
  assign _12004_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [10] : \MSYNC_1r1w.synth.nz.mem[706] [10];
  assign _12005_ = \bapg_rd.w_ptr_r [1] ? _12004_ : _12003_;
  assign _12006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [10] : \MSYNC_1r1w.synth.nz.mem[708] [10];
  assign _12007_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [10] : \MSYNC_1r1w.synth.nz.mem[710] [10];
  assign _12008_ = \bapg_rd.w_ptr_r [1] ? _12007_ : _12006_;
  assign _12009_ = \bapg_rd.w_ptr_r [2] ? _12008_ : _12005_;
  assign _12010_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [10] : \MSYNC_1r1w.synth.nz.mem[712] [10];
  assign _12011_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [10] : \MSYNC_1r1w.synth.nz.mem[714] [10];
  assign _12012_ = \bapg_rd.w_ptr_r [1] ? _12011_ : _12010_;
  assign _12013_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [10] : \MSYNC_1r1w.synth.nz.mem[716] [10];
  assign _12014_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [10] : \MSYNC_1r1w.synth.nz.mem[718] [10];
  assign _12015_ = \bapg_rd.w_ptr_r [1] ? _12014_ : _12013_;
  assign _12016_ = \bapg_rd.w_ptr_r [2] ? _12015_ : _12012_;
  assign _12017_ = \bapg_rd.w_ptr_r [3] ? _12016_ : _12009_;
  assign _12018_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [10] : \MSYNC_1r1w.synth.nz.mem[720] [10];
  assign _12019_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [10] : \MSYNC_1r1w.synth.nz.mem[722] [10];
  assign _12020_ = \bapg_rd.w_ptr_r [1] ? _12019_ : _12018_;
  assign _12021_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [10] : \MSYNC_1r1w.synth.nz.mem[724] [10];
  assign _12022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [10] : \MSYNC_1r1w.synth.nz.mem[726] [10];
  assign _12023_ = \bapg_rd.w_ptr_r [1] ? _12022_ : _12021_;
  assign _12024_ = \bapg_rd.w_ptr_r [2] ? _12023_ : _12020_;
  assign _12025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [10] : \MSYNC_1r1w.synth.nz.mem[728] [10];
  assign _12026_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [10] : \MSYNC_1r1w.synth.nz.mem[730] [10];
  assign _12027_ = \bapg_rd.w_ptr_r [1] ? _12026_ : _12025_;
  assign _12028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [10] : \MSYNC_1r1w.synth.nz.mem[732] [10];
  assign _12029_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [10] : \MSYNC_1r1w.synth.nz.mem[734] [10];
  assign _12030_ = \bapg_rd.w_ptr_r [1] ? _12029_ : _12028_;
  assign _12031_ = \bapg_rd.w_ptr_r [2] ? _12030_ : _12027_;
  assign _12032_ = \bapg_rd.w_ptr_r [3] ? _12031_ : _12024_;
  assign _12033_ = \bapg_rd.w_ptr_r [4] ? _12032_ : _12017_;
  assign _12034_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [10] : \MSYNC_1r1w.synth.nz.mem[736] [10];
  assign _12035_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [10] : \MSYNC_1r1w.synth.nz.mem[738] [10];
  assign _12036_ = \bapg_rd.w_ptr_r [1] ? _12035_ : _12034_;
  assign _12037_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [10] : \MSYNC_1r1w.synth.nz.mem[740] [10];
  assign _12038_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [10] : \MSYNC_1r1w.synth.nz.mem[742] [10];
  assign _12039_ = \bapg_rd.w_ptr_r [1] ? _12038_ : _12037_;
  assign _12040_ = \bapg_rd.w_ptr_r [2] ? _12039_ : _12036_;
  assign _12041_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [10] : \MSYNC_1r1w.synth.nz.mem[744] [10];
  assign _12042_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [10] : \MSYNC_1r1w.synth.nz.mem[746] [10];
  assign _12043_ = \bapg_rd.w_ptr_r [1] ? _12042_ : _12041_;
  assign _12044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [10] : \MSYNC_1r1w.synth.nz.mem[748] [10];
  assign _12045_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [10] : \MSYNC_1r1w.synth.nz.mem[750] [10];
  assign _12046_ = \bapg_rd.w_ptr_r [1] ? _12045_ : _12044_;
  assign _12047_ = \bapg_rd.w_ptr_r [2] ? _12046_ : _12043_;
  assign _12048_ = \bapg_rd.w_ptr_r [3] ? _12047_ : _12040_;
  assign _12049_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [10] : \MSYNC_1r1w.synth.nz.mem[752] [10];
  assign _12050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [10] : \MSYNC_1r1w.synth.nz.mem[754] [10];
  assign _12051_ = \bapg_rd.w_ptr_r [1] ? _12050_ : _12049_;
  assign _12052_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [10] : \MSYNC_1r1w.synth.nz.mem[756] [10];
  assign _12053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [10] : \MSYNC_1r1w.synth.nz.mem[758] [10];
  assign _12054_ = \bapg_rd.w_ptr_r [1] ? _12053_ : _12052_;
  assign _12055_ = \bapg_rd.w_ptr_r [2] ? _12054_ : _12051_;
  assign _12056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [10] : \MSYNC_1r1w.synth.nz.mem[760] [10];
  assign _12057_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [10] : \MSYNC_1r1w.synth.nz.mem[762] [10];
  assign _12058_ = \bapg_rd.w_ptr_r [1] ? _12057_ : _12056_;
  assign _12059_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [10] : \MSYNC_1r1w.synth.nz.mem[764] [10];
  assign _12060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [10] : \MSYNC_1r1w.synth.nz.mem[766] [10];
  assign _12061_ = \bapg_rd.w_ptr_r [1] ? _12060_ : _12059_;
  assign _12062_ = \bapg_rd.w_ptr_r [2] ? _12061_ : _12058_;
  assign _12063_ = \bapg_rd.w_ptr_r [3] ? _12062_ : _12055_;
  assign _12064_ = \bapg_rd.w_ptr_r [4] ? _12063_ : _12048_;
  assign _12065_ = \bapg_rd.w_ptr_r [5] ? _12064_ : _12033_;
  assign _12066_ = \bapg_rd.w_ptr_r [6] ? _12065_ : _12002_;
  assign _12067_ = \bapg_rd.w_ptr_r [7] ? _12066_ : _11939_;
  assign _12068_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [10] : \MSYNC_1r1w.synth.nz.mem[768] [10];
  assign _12069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [10] : \MSYNC_1r1w.synth.nz.mem[770] [10];
  assign _12070_ = \bapg_rd.w_ptr_r [1] ? _12069_ : _12068_;
  assign _12071_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [10] : \MSYNC_1r1w.synth.nz.mem[772] [10];
  assign _12072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [10] : \MSYNC_1r1w.synth.nz.mem[774] [10];
  assign _12073_ = \bapg_rd.w_ptr_r [1] ? _12072_ : _12071_;
  assign _12074_ = \bapg_rd.w_ptr_r [2] ? _12073_ : _12070_;
  assign _12075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [10] : \MSYNC_1r1w.synth.nz.mem[776] [10];
  assign _12076_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [10] : \MSYNC_1r1w.synth.nz.mem[778] [10];
  assign _12077_ = \bapg_rd.w_ptr_r [1] ? _12076_ : _12075_;
  assign _12078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [10] : \MSYNC_1r1w.synth.nz.mem[780] [10];
  assign _12079_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [10] : \MSYNC_1r1w.synth.nz.mem[782] [10];
  assign _12080_ = \bapg_rd.w_ptr_r [1] ? _12079_ : _12078_;
  assign _12081_ = \bapg_rd.w_ptr_r [2] ? _12080_ : _12077_;
  assign _12082_ = \bapg_rd.w_ptr_r [3] ? _12081_ : _12074_;
  assign _12083_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [10] : \MSYNC_1r1w.synth.nz.mem[784] [10];
  assign _12084_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [10] : \MSYNC_1r1w.synth.nz.mem[786] [10];
  assign _12085_ = \bapg_rd.w_ptr_r [1] ? _12084_ : _12083_;
  assign _12086_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [10] : \MSYNC_1r1w.synth.nz.mem[788] [10];
  assign _12087_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [10] : \MSYNC_1r1w.synth.nz.mem[790] [10];
  assign _12088_ = \bapg_rd.w_ptr_r [1] ? _12087_ : _12086_;
  assign _12089_ = \bapg_rd.w_ptr_r [2] ? _12088_ : _12085_;
  assign _12090_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [10] : \MSYNC_1r1w.synth.nz.mem[792] [10];
  assign _12091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [10] : \MSYNC_1r1w.synth.nz.mem[794] [10];
  assign _12092_ = \bapg_rd.w_ptr_r [1] ? _12091_ : _12090_;
  assign _12093_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [10] : \MSYNC_1r1w.synth.nz.mem[796] [10];
  assign _12094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [10] : \MSYNC_1r1w.synth.nz.mem[798] [10];
  assign _12095_ = \bapg_rd.w_ptr_r [1] ? _12094_ : _12093_;
  assign _12096_ = \bapg_rd.w_ptr_r [2] ? _12095_ : _12092_;
  assign _12097_ = \bapg_rd.w_ptr_r [3] ? _12096_ : _12089_;
  assign _12098_ = \bapg_rd.w_ptr_r [4] ? _12097_ : _12082_;
  assign _12099_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [10] : \MSYNC_1r1w.synth.nz.mem[800] [10];
  assign _12100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [10] : \MSYNC_1r1w.synth.nz.mem[802] [10];
  assign _12101_ = \bapg_rd.w_ptr_r [1] ? _12100_ : _12099_;
  assign _12102_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [10] : \MSYNC_1r1w.synth.nz.mem[804] [10];
  assign _12103_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [10] : \MSYNC_1r1w.synth.nz.mem[806] [10];
  assign _12104_ = \bapg_rd.w_ptr_r [1] ? _12103_ : _12102_;
  assign _12105_ = \bapg_rd.w_ptr_r [2] ? _12104_ : _12101_;
  assign _12106_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [10] : \MSYNC_1r1w.synth.nz.mem[808] [10];
  assign _12107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [10] : \MSYNC_1r1w.synth.nz.mem[810] [10];
  assign _12108_ = \bapg_rd.w_ptr_r [1] ? _12107_ : _12106_;
  assign _12109_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [10] : \MSYNC_1r1w.synth.nz.mem[812] [10];
  assign _12110_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [10] : \MSYNC_1r1w.synth.nz.mem[814] [10];
  assign _12111_ = \bapg_rd.w_ptr_r [1] ? _12110_ : _12109_;
  assign _12112_ = \bapg_rd.w_ptr_r [2] ? _12111_ : _12108_;
  assign _12113_ = \bapg_rd.w_ptr_r [3] ? _12112_ : _12105_;
  assign _12114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [10] : \MSYNC_1r1w.synth.nz.mem[816] [10];
  assign _12115_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [10] : \MSYNC_1r1w.synth.nz.mem[818] [10];
  assign _12116_ = \bapg_rd.w_ptr_r [1] ? _12115_ : _12114_;
  assign _12117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [10] : \MSYNC_1r1w.synth.nz.mem[820] [10];
  assign _12118_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [10] : \MSYNC_1r1w.synth.nz.mem[822] [10];
  assign _12119_ = \bapg_rd.w_ptr_r [1] ? _12118_ : _12117_;
  assign _12120_ = \bapg_rd.w_ptr_r [2] ? _12119_ : _12116_;
  assign _12121_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [10] : \MSYNC_1r1w.synth.nz.mem[824] [10];
  assign _12122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [10] : \MSYNC_1r1w.synth.nz.mem[826] [10];
  assign _12123_ = \bapg_rd.w_ptr_r [1] ? _12122_ : _12121_;
  assign _12124_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [10] : \MSYNC_1r1w.synth.nz.mem[828] [10];
  assign _12125_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [10] : \MSYNC_1r1w.synth.nz.mem[830] [10];
  assign _12126_ = \bapg_rd.w_ptr_r [1] ? _12125_ : _12124_;
  assign _12127_ = \bapg_rd.w_ptr_r [2] ? _12126_ : _12123_;
  assign _12128_ = \bapg_rd.w_ptr_r [3] ? _12127_ : _12120_;
  assign _12129_ = \bapg_rd.w_ptr_r [4] ? _12128_ : _12113_;
  assign _12130_ = \bapg_rd.w_ptr_r [5] ? _12129_ : _12098_;
  assign _12131_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [10] : \MSYNC_1r1w.synth.nz.mem[832] [10];
  assign _12132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [10] : \MSYNC_1r1w.synth.nz.mem[834] [10];
  assign _12133_ = \bapg_rd.w_ptr_r [1] ? _12132_ : _12131_;
  assign _12134_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [10] : \MSYNC_1r1w.synth.nz.mem[836] [10];
  assign _12135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [10] : \MSYNC_1r1w.synth.nz.mem[838] [10];
  assign _12136_ = \bapg_rd.w_ptr_r [1] ? _12135_ : _12134_;
  assign _12137_ = \bapg_rd.w_ptr_r [2] ? _12136_ : _12133_;
  assign _12138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [10] : \MSYNC_1r1w.synth.nz.mem[840] [10];
  assign _12139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [10] : \MSYNC_1r1w.synth.nz.mem[842] [10];
  assign _12140_ = \bapg_rd.w_ptr_r [1] ? _12139_ : _12138_;
  assign _12141_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [10] : \MSYNC_1r1w.synth.nz.mem[844] [10];
  assign _12142_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [10] : \MSYNC_1r1w.synth.nz.mem[846] [10];
  assign _12143_ = \bapg_rd.w_ptr_r [1] ? _12142_ : _12141_;
  assign _12144_ = \bapg_rd.w_ptr_r [2] ? _12143_ : _12140_;
  assign _12145_ = \bapg_rd.w_ptr_r [3] ? _12144_ : _12137_;
  assign _12146_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [10] : \MSYNC_1r1w.synth.nz.mem[848] [10];
  assign _12147_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [10] : \MSYNC_1r1w.synth.nz.mem[850] [10];
  assign _12148_ = \bapg_rd.w_ptr_r [1] ? _12147_ : _12146_;
  assign _12149_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [10] : \MSYNC_1r1w.synth.nz.mem[852] [10];
  assign _12150_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [10] : \MSYNC_1r1w.synth.nz.mem[854] [10];
  assign _12151_ = \bapg_rd.w_ptr_r [1] ? _12150_ : _12149_;
  assign _12152_ = \bapg_rd.w_ptr_r [2] ? _12151_ : _12148_;
  assign _12153_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [10] : \MSYNC_1r1w.synth.nz.mem[856] [10];
  assign _12154_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [10] : \MSYNC_1r1w.synth.nz.mem[858] [10];
  assign _12155_ = \bapg_rd.w_ptr_r [1] ? _12154_ : _12153_;
  assign _12156_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [10] : \MSYNC_1r1w.synth.nz.mem[860] [10];
  assign _12157_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [10] : \MSYNC_1r1w.synth.nz.mem[862] [10];
  assign _12158_ = \bapg_rd.w_ptr_r [1] ? _12157_ : _12156_;
  assign _12159_ = \bapg_rd.w_ptr_r [2] ? _12158_ : _12155_;
  assign _12160_ = \bapg_rd.w_ptr_r [3] ? _12159_ : _12152_;
  assign _12161_ = \bapg_rd.w_ptr_r [4] ? _12160_ : _12145_;
  assign _12162_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [10] : \MSYNC_1r1w.synth.nz.mem[864] [10];
  assign _12163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [10] : \MSYNC_1r1w.synth.nz.mem[866] [10];
  assign _12164_ = \bapg_rd.w_ptr_r [1] ? _12163_ : _12162_;
  assign _12165_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [10] : \MSYNC_1r1w.synth.nz.mem[868] [10];
  assign _12166_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [10] : \MSYNC_1r1w.synth.nz.mem[870] [10];
  assign _12167_ = \bapg_rd.w_ptr_r [1] ? _12166_ : _12165_;
  assign _12168_ = \bapg_rd.w_ptr_r [2] ? _12167_ : _12164_;
  assign _12169_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [10] : \MSYNC_1r1w.synth.nz.mem[872] [10];
  assign _12170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [10] : \MSYNC_1r1w.synth.nz.mem[874] [10];
  assign _12171_ = \bapg_rd.w_ptr_r [1] ? _12170_ : _12169_;
  assign _12172_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [10] : \MSYNC_1r1w.synth.nz.mem[876] [10];
  assign _12173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [10] : \MSYNC_1r1w.synth.nz.mem[878] [10];
  assign _12174_ = \bapg_rd.w_ptr_r [1] ? _12173_ : _12172_;
  assign _12175_ = \bapg_rd.w_ptr_r [2] ? _12174_ : _12171_;
  assign _12176_ = \bapg_rd.w_ptr_r [3] ? _12175_ : _12168_;
  assign _12177_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [10] : \MSYNC_1r1w.synth.nz.mem[880] [10];
  assign _12178_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [10] : \MSYNC_1r1w.synth.nz.mem[882] [10];
  assign _12179_ = \bapg_rd.w_ptr_r [1] ? _12178_ : _12177_;
  assign _12180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [10] : \MSYNC_1r1w.synth.nz.mem[884] [10];
  assign _12181_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [10] : \MSYNC_1r1w.synth.nz.mem[886] [10];
  assign _12182_ = \bapg_rd.w_ptr_r [1] ? _12181_ : _12180_;
  assign _12183_ = \bapg_rd.w_ptr_r [2] ? _12182_ : _12179_;
  assign _12184_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [10] : \MSYNC_1r1w.synth.nz.mem[888] [10];
  assign _12185_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [10] : \MSYNC_1r1w.synth.nz.mem[890] [10];
  assign _12186_ = \bapg_rd.w_ptr_r [1] ? _12185_ : _12184_;
  assign _12187_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [10] : \MSYNC_1r1w.synth.nz.mem[892] [10];
  assign _12188_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [10] : \MSYNC_1r1w.synth.nz.mem[894] [10];
  assign _12189_ = \bapg_rd.w_ptr_r [1] ? _12188_ : _12187_;
  assign _12190_ = \bapg_rd.w_ptr_r [2] ? _12189_ : _12186_;
  assign _12191_ = \bapg_rd.w_ptr_r [3] ? _12190_ : _12183_;
  assign _12192_ = \bapg_rd.w_ptr_r [4] ? _12191_ : _12176_;
  assign _12193_ = \bapg_rd.w_ptr_r [5] ? _12192_ : _12161_;
  assign _12194_ = \bapg_rd.w_ptr_r [6] ? _12193_ : _12130_;
  assign _12195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [10] : \MSYNC_1r1w.synth.nz.mem[896] [10];
  assign _12196_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [10] : \MSYNC_1r1w.synth.nz.mem[898] [10];
  assign _12197_ = \bapg_rd.w_ptr_r [1] ? _12196_ : _12195_;
  assign _12198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [10] : \MSYNC_1r1w.synth.nz.mem[900] [10];
  assign _12199_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [10] : \MSYNC_1r1w.synth.nz.mem[902] [10];
  assign _12200_ = \bapg_rd.w_ptr_r [1] ? _12199_ : _12198_;
  assign _12201_ = \bapg_rd.w_ptr_r [2] ? _12200_ : _12197_;
  assign _12202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [10] : \MSYNC_1r1w.synth.nz.mem[904] [10];
  assign _12203_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [10] : \MSYNC_1r1w.synth.nz.mem[906] [10];
  assign _12204_ = \bapg_rd.w_ptr_r [1] ? _12203_ : _12202_;
  assign _12205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [10] : \MSYNC_1r1w.synth.nz.mem[908] [10];
  assign _12206_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [10] : \MSYNC_1r1w.synth.nz.mem[910] [10];
  assign _12207_ = \bapg_rd.w_ptr_r [1] ? _12206_ : _12205_;
  assign _12208_ = \bapg_rd.w_ptr_r [2] ? _12207_ : _12204_;
  assign _12209_ = \bapg_rd.w_ptr_r [3] ? _12208_ : _12201_;
  assign _12210_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [10] : \MSYNC_1r1w.synth.nz.mem[912] [10];
  assign _12211_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [10] : \MSYNC_1r1w.synth.nz.mem[914] [10];
  assign _12212_ = \bapg_rd.w_ptr_r [1] ? _12211_ : _12210_;
  assign _12213_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [10] : \MSYNC_1r1w.synth.nz.mem[916] [10];
  assign _12214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [10] : \MSYNC_1r1w.synth.nz.mem[918] [10];
  assign _12215_ = \bapg_rd.w_ptr_r [1] ? _12214_ : _12213_;
  assign _12216_ = \bapg_rd.w_ptr_r [2] ? _12215_ : _12212_;
  assign _12217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [10] : \MSYNC_1r1w.synth.nz.mem[920] [10];
  assign _12218_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [10] : \MSYNC_1r1w.synth.nz.mem[922] [10];
  assign _12219_ = \bapg_rd.w_ptr_r [1] ? _12218_ : _12217_;
  assign _12220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [10] : \MSYNC_1r1w.synth.nz.mem[924] [10];
  assign _12221_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [10] : \MSYNC_1r1w.synth.nz.mem[926] [10];
  assign _12222_ = \bapg_rd.w_ptr_r [1] ? _12221_ : _12220_;
  assign _12223_ = \bapg_rd.w_ptr_r [2] ? _12222_ : _12219_;
  assign _12224_ = \bapg_rd.w_ptr_r [3] ? _12223_ : _12216_;
  assign _12225_ = \bapg_rd.w_ptr_r [4] ? _12224_ : _12209_;
  assign _12226_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [10] : \MSYNC_1r1w.synth.nz.mem[928] [10];
  assign _12227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [10] : \MSYNC_1r1w.synth.nz.mem[930] [10];
  assign _12228_ = \bapg_rd.w_ptr_r [1] ? _12227_ : _12226_;
  assign _12229_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [10] : \MSYNC_1r1w.synth.nz.mem[932] [10];
  assign _12230_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [10] : \MSYNC_1r1w.synth.nz.mem[934] [10];
  assign _12231_ = \bapg_rd.w_ptr_r [1] ? _12230_ : _12229_;
  assign _12232_ = \bapg_rd.w_ptr_r [2] ? _12231_ : _12228_;
  assign _12233_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [10] : \MSYNC_1r1w.synth.nz.mem[936] [10];
  assign _12234_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [10] : \MSYNC_1r1w.synth.nz.mem[938] [10];
  assign _12235_ = \bapg_rd.w_ptr_r [1] ? _12234_ : _12233_;
  assign _12236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [10] : \MSYNC_1r1w.synth.nz.mem[940] [10];
  assign _12237_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [10] : \MSYNC_1r1w.synth.nz.mem[942] [10];
  assign _12238_ = \bapg_rd.w_ptr_r [1] ? _12237_ : _12236_;
  assign _12239_ = \bapg_rd.w_ptr_r [2] ? _12238_ : _12235_;
  assign _12240_ = \bapg_rd.w_ptr_r [3] ? _12239_ : _12232_;
  assign _12241_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [10] : \MSYNC_1r1w.synth.nz.mem[944] [10];
  assign _12242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [10] : \MSYNC_1r1w.synth.nz.mem[946] [10];
  assign _12243_ = \bapg_rd.w_ptr_r [1] ? _12242_ : _12241_;
  assign _12244_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [10] : \MSYNC_1r1w.synth.nz.mem[948] [10];
  assign _12245_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [10] : \MSYNC_1r1w.synth.nz.mem[950] [10];
  assign _12246_ = \bapg_rd.w_ptr_r [1] ? _12245_ : _12244_;
  assign _12247_ = \bapg_rd.w_ptr_r [2] ? _12246_ : _12243_;
  assign _12248_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [10] : \MSYNC_1r1w.synth.nz.mem[952] [10];
  assign _12249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [10] : \MSYNC_1r1w.synth.nz.mem[954] [10];
  assign _12250_ = \bapg_rd.w_ptr_r [1] ? _12249_ : _12248_;
  assign _12251_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [10] : \MSYNC_1r1w.synth.nz.mem[956] [10];
  assign _12252_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [10] : \MSYNC_1r1w.synth.nz.mem[958] [10];
  assign _12253_ = \bapg_rd.w_ptr_r [1] ? _12252_ : _12251_;
  assign _12254_ = \bapg_rd.w_ptr_r [2] ? _12253_ : _12250_;
  assign _12255_ = \bapg_rd.w_ptr_r [3] ? _12254_ : _12247_;
  assign _12256_ = \bapg_rd.w_ptr_r [4] ? _12255_ : _12240_;
  assign _12257_ = \bapg_rd.w_ptr_r [5] ? _12256_ : _12225_;
  assign _12258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [10] : \MSYNC_1r1w.synth.nz.mem[960] [10];
  assign _12259_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [10] : \MSYNC_1r1w.synth.nz.mem[962] [10];
  assign _12260_ = \bapg_rd.w_ptr_r [1] ? _12259_ : _12258_;
  assign _12261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [10] : \MSYNC_1r1w.synth.nz.mem[964] [10];
  assign _12262_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [10] : \MSYNC_1r1w.synth.nz.mem[966] [10];
  assign _12263_ = \bapg_rd.w_ptr_r [1] ? _12262_ : _12261_;
  assign _12264_ = \bapg_rd.w_ptr_r [2] ? _12263_ : _12260_;
  assign _12265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [10] : \MSYNC_1r1w.synth.nz.mem[968] [10];
  assign _12266_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [10] : \MSYNC_1r1w.synth.nz.mem[970] [10];
  assign _12267_ = \bapg_rd.w_ptr_r [1] ? _12266_ : _12265_;
  assign _12268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [10] : \MSYNC_1r1w.synth.nz.mem[972] [10];
  assign _12269_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [10] : \MSYNC_1r1w.synth.nz.mem[974] [10];
  assign _12270_ = \bapg_rd.w_ptr_r [1] ? _12269_ : _12268_;
  assign _12271_ = \bapg_rd.w_ptr_r [2] ? _12270_ : _12267_;
  assign _12272_ = \bapg_rd.w_ptr_r [3] ? _12271_ : _12264_;
  assign _12273_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [10] : \MSYNC_1r1w.synth.nz.mem[976] [10];
  assign _12274_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [10] : \MSYNC_1r1w.synth.nz.mem[978] [10];
  assign _12275_ = \bapg_rd.w_ptr_r [1] ? _12274_ : _12273_;
  assign _12276_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [10] : \MSYNC_1r1w.synth.nz.mem[980] [10];
  assign _12277_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [10] : \MSYNC_1r1w.synth.nz.mem[982] [10];
  assign _12278_ = \bapg_rd.w_ptr_r [1] ? _12277_ : _12276_;
  assign _12279_ = \bapg_rd.w_ptr_r [2] ? _12278_ : _12275_;
  assign _12280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [10] : \MSYNC_1r1w.synth.nz.mem[984] [10];
  assign _12281_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [10] : \MSYNC_1r1w.synth.nz.mem[986] [10];
  assign _12282_ = \bapg_rd.w_ptr_r [1] ? _12281_ : _12280_;
  assign _12283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [10] : \MSYNC_1r1w.synth.nz.mem[988] [10];
  assign _12284_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [10] : \MSYNC_1r1w.synth.nz.mem[990] [10];
  assign _12285_ = \bapg_rd.w_ptr_r [1] ? _12284_ : _12283_;
  assign _12286_ = \bapg_rd.w_ptr_r [2] ? _12285_ : _12282_;
  assign _12287_ = \bapg_rd.w_ptr_r [3] ? _12286_ : _12279_;
  assign _12288_ = \bapg_rd.w_ptr_r [4] ? _12287_ : _12272_;
  assign _12289_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [10] : \MSYNC_1r1w.synth.nz.mem[992] [10];
  assign _12290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [10] : \MSYNC_1r1w.synth.nz.mem[994] [10];
  assign _12291_ = \bapg_rd.w_ptr_r [1] ? _12290_ : _12289_;
  assign _12292_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [10] : \MSYNC_1r1w.synth.nz.mem[996] [10];
  assign _12293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [10] : \MSYNC_1r1w.synth.nz.mem[998] [10];
  assign _12294_ = \bapg_rd.w_ptr_r [1] ? _12293_ : _12292_;
  assign _12295_ = \bapg_rd.w_ptr_r [2] ? _12294_ : _12291_;
  assign _12296_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [10] : \MSYNC_1r1w.synth.nz.mem[1000] [10];
  assign _12297_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [10] : \MSYNC_1r1w.synth.nz.mem[1002] [10];
  assign _12298_ = \bapg_rd.w_ptr_r [1] ? _12297_ : _12296_;
  assign _12299_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [10] : \MSYNC_1r1w.synth.nz.mem[1004] [10];
  assign _12300_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [10] : \MSYNC_1r1w.synth.nz.mem[1006] [10];
  assign _12301_ = \bapg_rd.w_ptr_r [1] ? _12300_ : _12299_;
  assign _12302_ = \bapg_rd.w_ptr_r [2] ? _12301_ : _12298_;
  assign _12303_ = \bapg_rd.w_ptr_r [3] ? _12302_ : _12295_;
  assign _12304_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [10] : \MSYNC_1r1w.synth.nz.mem[1008] [10];
  assign _12305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [10] : \MSYNC_1r1w.synth.nz.mem[1010] [10];
  assign _12306_ = \bapg_rd.w_ptr_r [1] ? _12305_ : _12304_;
  assign _12307_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [10] : \MSYNC_1r1w.synth.nz.mem[1012] [10];
  assign _12308_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [10] : \MSYNC_1r1w.synth.nz.mem[1014] [10];
  assign _12309_ = \bapg_rd.w_ptr_r [1] ? _12308_ : _12307_;
  assign _12310_ = \bapg_rd.w_ptr_r [2] ? _12309_ : _12306_;
  assign _12311_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [10] : \MSYNC_1r1w.synth.nz.mem[1016] [10];
  assign _12312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [10] : \MSYNC_1r1w.synth.nz.mem[1018] [10];
  assign _12313_ = \bapg_rd.w_ptr_r [1] ? _12312_ : _12311_;
  assign _12314_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [10] : \MSYNC_1r1w.synth.nz.mem[1020] [10];
  assign _12315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [10] : \MSYNC_1r1w.synth.nz.mem[1022] [10];
  assign _12316_ = \bapg_rd.w_ptr_r [1] ? _12315_ : _12314_;
  assign _12317_ = \bapg_rd.w_ptr_r [2] ? _12316_ : _12313_;
  assign _12318_ = \bapg_rd.w_ptr_r [3] ? _12317_ : _12310_;
  assign _12319_ = \bapg_rd.w_ptr_r [4] ? _12318_ : _12303_;
  assign _12320_ = \bapg_rd.w_ptr_r [5] ? _12319_ : _12288_;
  assign _12321_ = \bapg_rd.w_ptr_r [6] ? _12320_ : _12257_;
  assign _12322_ = \bapg_rd.w_ptr_r [7] ? _12321_ : _12194_;
  assign _12323_ = \bapg_rd.w_ptr_r [8] ? _12322_ : _12067_;
  assign r_data_o[10] = \bapg_rd.w_ptr_r [9] ? _12323_ : _11812_;
  assign _12324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [11] : \MSYNC_1r1w.synth.nz.mem[0] [11];
  assign _12325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [11] : \MSYNC_1r1w.synth.nz.mem[2] [11];
  assign _12326_ = \bapg_rd.w_ptr_r [1] ? _12325_ : _12324_;
  assign _12327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [11] : \MSYNC_1r1w.synth.nz.mem[4] [11];
  assign _12328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [11] : \MSYNC_1r1w.synth.nz.mem[6] [11];
  assign _12329_ = \bapg_rd.w_ptr_r [1] ? _12328_ : _12327_;
  assign _12330_ = \bapg_rd.w_ptr_r [2] ? _12329_ : _12326_;
  assign _12331_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [11] : \MSYNC_1r1w.synth.nz.mem[8] [11];
  assign _12332_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [11] : \MSYNC_1r1w.synth.nz.mem[10] [11];
  assign _12333_ = \bapg_rd.w_ptr_r [1] ? _12332_ : _12331_;
  assign _12334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [11] : \MSYNC_1r1w.synth.nz.mem[12] [11];
  assign _12335_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [11] : \MSYNC_1r1w.synth.nz.mem[14] [11];
  assign _12336_ = \bapg_rd.w_ptr_r [1] ? _12335_ : _12334_;
  assign _12337_ = \bapg_rd.w_ptr_r [2] ? _12336_ : _12333_;
  assign _12338_ = \bapg_rd.w_ptr_r [3] ? _12337_ : _12330_;
  assign _12339_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [11] : \MSYNC_1r1w.synth.nz.mem[16] [11];
  assign _12340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [11] : \MSYNC_1r1w.synth.nz.mem[18] [11];
  assign _12341_ = \bapg_rd.w_ptr_r [1] ? _12340_ : _12339_;
  assign _12342_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [11] : \MSYNC_1r1w.synth.nz.mem[20] [11];
  assign _12343_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [11] : \MSYNC_1r1w.synth.nz.mem[22] [11];
  assign _12344_ = \bapg_rd.w_ptr_r [1] ? _12343_ : _12342_;
  assign _12345_ = \bapg_rd.w_ptr_r [2] ? _12344_ : _12341_;
  assign _12346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [11] : \MSYNC_1r1w.synth.nz.mem[24] [11];
  assign _12347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [11] : \MSYNC_1r1w.synth.nz.mem[26] [11];
  assign _12348_ = \bapg_rd.w_ptr_r [1] ? _12347_ : _12346_;
  assign _12349_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [11] : \MSYNC_1r1w.synth.nz.mem[28] [11];
  assign _12350_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [11] : \MSYNC_1r1w.synth.nz.mem[30] [11];
  assign _12351_ = \bapg_rd.w_ptr_r [1] ? _12350_ : _12349_;
  assign _12352_ = \bapg_rd.w_ptr_r [2] ? _12351_ : _12348_;
  assign _12353_ = \bapg_rd.w_ptr_r [3] ? _12352_ : _12345_;
  assign _12354_ = \bapg_rd.w_ptr_r [4] ? _12353_ : _12338_;
  assign _12355_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [11] : \MSYNC_1r1w.synth.nz.mem[32] [11];
  assign _12356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [11] : \MSYNC_1r1w.synth.nz.mem[34] [11];
  assign _12357_ = \bapg_rd.w_ptr_r [1] ? _12356_ : _12355_;
  assign _12358_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [11] : \MSYNC_1r1w.synth.nz.mem[36] [11];
  assign _12359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [11] : \MSYNC_1r1w.synth.nz.mem[38] [11];
  assign _12360_ = \bapg_rd.w_ptr_r [1] ? _12359_ : _12358_;
  assign _12361_ = \bapg_rd.w_ptr_r [2] ? _12360_ : _12357_;
  assign _12362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [11] : \MSYNC_1r1w.synth.nz.mem[40] [11];
  assign _12363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [11] : \MSYNC_1r1w.synth.nz.mem[42] [11];
  assign _12364_ = \bapg_rd.w_ptr_r [1] ? _12363_ : _12362_;
  assign _12365_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [11] : \MSYNC_1r1w.synth.nz.mem[44] [11];
  assign _12366_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [11] : \MSYNC_1r1w.synth.nz.mem[46] [11];
  assign _12367_ = \bapg_rd.w_ptr_r [1] ? _12366_ : _12365_;
  assign _12368_ = \bapg_rd.w_ptr_r [2] ? _12367_ : _12364_;
  assign _12369_ = \bapg_rd.w_ptr_r [3] ? _12368_ : _12361_;
  assign _12370_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [11] : \MSYNC_1r1w.synth.nz.mem[48] [11];
  assign _12371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [11] : \MSYNC_1r1w.synth.nz.mem[50] [11];
  assign _12372_ = \bapg_rd.w_ptr_r [1] ? _12371_ : _12370_;
  assign _12373_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [11] : \MSYNC_1r1w.synth.nz.mem[52] [11];
  assign _12374_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [11] : \MSYNC_1r1w.synth.nz.mem[54] [11];
  assign _12375_ = \bapg_rd.w_ptr_r [1] ? _12374_ : _12373_;
  assign _12376_ = \bapg_rd.w_ptr_r [2] ? _12375_ : _12372_;
  assign _12377_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [11] : \MSYNC_1r1w.synth.nz.mem[56] [11];
  assign _12378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [11] : \MSYNC_1r1w.synth.nz.mem[58] [11];
  assign _12379_ = \bapg_rd.w_ptr_r [1] ? _12378_ : _12377_;
  assign _12380_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [11] : \MSYNC_1r1w.synth.nz.mem[60] [11];
  assign _12381_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [11] : \MSYNC_1r1w.synth.nz.mem[62] [11];
  assign _12382_ = \bapg_rd.w_ptr_r [1] ? _12381_ : _12380_;
  assign _12383_ = \bapg_rd.w_ptr_r [2] ? _12382_ : _12379_;
  assign _12384_ = \bapg_rd.w_ptr_r [3] ? _12383_ : _12376_;
  assign _12385_ = \bapg_rd.w_ptr_r [4] ? _12384_ : _12369_;
  assign _12386_ = \bapg_rd.w_ptr_r [5] ? _12385_ : _12354_;
  assign _12387_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [11] : \MSYNC_1r1w.synth.nz.mem[64] [11];
  assign _12388_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [11] : \MSYNC_1r1w.synth.nz.mem[66] [11];
  assign _12389_ = \bapg_rd.w_ptr_r [1] ? _12388_ : _12387_;
  assign _12390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [11] : \MSYNC_1r1w.synth.nz.mem[68] [11];
  assign _12391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [11] : \MSYNC_1r1w.synth.nz.mem[70] [11];
  assign _12392_ = \bapg_rd.w_ptr_r [1] ? _12391_ : _12390_;
  assign _12393_ = \bapg_rd.w_ptr_r [2] ? _12392_ : _12389_;
  assign _12394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [11] : \MSYNC_1r1w.synth.nz.mem[72] [11];
  assign _12395_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [11] : \MSYNC_1r1w.synth.nz.mem[74] [11];
  assign _12396_ = \bapg_rd.w_ptr_r [1] ? _12395_ : _12394_;
  assign _12397_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [11] : \MSYNC_1r1w.synth.nz.mem[76] [11];
  assign _12398_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [11] : \MSYNC_1r1w.synth.nz.mem[78] [11];
  assign _12399_ = \bapg_rd.w_ptr_r [1] ? _12398_ : _12397_;
  assign _12400_ = \bapg_rd.w_ptr_r [2] ? _12399_ : _12396_;
  assign _12401_ = \bapg_rd.w_ptr_r [3] ? _12400_ : _12393_;
  assign _12402_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [11] : \MSYNC_1r1w.synth.nz.mem[80] [11];
  assign _12403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [11] : \MSYNC_1r1w.synth.nz.mem[82] [11];
  assign _12404_ = \bapg_rd.w_ptr_r [1] ? _12403_ : _12402_;
  assign _12405_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [11] : \MSYNC_1r1w.synth.nz.mem[84] [11];
  assign _12406_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [11] : \MSYNC_1r1w.synth.nz.mem[86] [11];
  assign _12407_ = \bapg_rd.w_ptr_r [1] ? _12406_ : _12405_;
  assign _12408_ = \bapg_rd.w_ptr_r [2] ? _12407_ : _12404_;
  assign _12409_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [11] : \MSYNC_1r1w.synth.nz.mem[88] [11];
  assign _12410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [11] : \MSYNC_1r1w.synth.nz.mem[90] [11];
  assign _12411_ = \bapg_rd.w_ptr_r [1] ? _12410_ : _12409_;
  assign _12412_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [11] : \MSYNC_1r1w.synth.nz.mem[92] [11];
  assign _12413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [11] : \MSYNC_1r1w.synth.nz.mem[94] [11];
  assign _12414_ = \bapg_rd.w_ptr_r [1] ? _12413_ : _12412_;
  assign _12415_ = \bapg_rd.w_ptr_r [2] ? _12414_ : _12411_;
  assign _12416_ = \bapg_rd.w_ptr_r [3] ? _12415_ : _12408_;
  assign _12417_ = \bapg_rd.w_ptr_r [4] ? _12416_ : _12401_;
  assign _12418_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [11] : \MSYNC_1r1w.synth.nz.mem[96] [11];
  assign _12419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [11] : \MSYNC_1r1w.synth.nz.mem[98] [11];
  assign _12420_ = \bapg_rd.w_ptr_r [1] ? _12419_ : _12418_;
  assign _12421_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [11] : \MSYNC_1r1w.synth.nz.mem[100] [11];
  assign _12422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [11] : \MSYNC_1r1w.synth.nz.mem[102] [11];
  assign _12423_ = \bapg_rd.w_ptr_r [1] ? _12422_ : _12421_;
  assign _12424_ = \bapg_rd.w_ptr_r [2] ? _12423_ : _12420_;
  assign _12425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [11] : \MSYNC_1r1w.synth.nz.mem[104] [11];
  assign _12426_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [11] : \MSYNC_1r1w.synth.nz.mem[106] [11];
  assign _12427_ = \bapg_rd.w_ptr_r [1] ? _12426_ : _12425_;
  assign _12428_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [11] : \MSYNC_1r1w.synth.nz.mem[108] [11];
  assign _12429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [11] : \MSYNC_1r1w.synth.nz.mem[110] [11];
  assign _12430_ = \bapg_rd.w_ptr_r [1] ? _12429_ : _12428_;
  assign _12431_ = \bapg_rd.w_ptr_r [2] ? _12430_ : _12427_;
  assign _12432_ = \bapg_rd.w_ptr_r [3] ? _12431_ : _12424_;
  assign _12433_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [11] : \MSYNC_1r1w.synth.nz.mem[112] [11];
  assign _12434_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [11] : \MSYNC_1r1w.synth.nz.mem[114] [11];
  assign _12435_ = \bapg_rd.w_ptr_r [1] ? _12434_ : _12433_;
  assign _12436_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [11] : \MSYNC_1r1w.synth.nz.mem[116] [11];
  assign _12437_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [11] : \MSYNC_1r1w.synth.nz.mem[118] [11];
  assign _12438_ = \bapg_rd.w_ptr_r [1] ? _12437_ : _12436_;
  assign _12439_ = \bapg_rd.w_ptr_r [2] ? _12438_ : _12435_;
  assign _12440_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [11] : \MSYNC_1r1w.synth.nz.mem[120] [11];
  assign _12441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [11] : \MSYNC_1r1w.synth.nz.mem[122] [11];
  assign _12442_ = \bapg_rd.w_ptr_r [1] ? _12441_ : _12440_;
  assign _12443_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [11] : \MSYNC_1r1w.synth.nz.mem[124] [11];
  assign _12444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [11] : \MSYNC_1r1w.synth.nz.mem[126] [11];
  assign _12445_ = \bapg_rd.w_ptr_r [1] ? _12444_ : _12443_;
  assign _12446_ = \bapg_rd.w_ptr_r [2] ? _12445_ : _12442_;
  assign _12447_ = \bapg_rd.w_ptr_r [3] ? _12446_ : _12439_;
  assign _12448_ = \bapg_rd.w_ptr_r [4] ? _12447_ : _12432_;
  assign _12449_ = \bapg_rd.w_ptr_r [5] ? _12448_ : _12417_;
  assign _12450_ = \bapg_rd.w_ptr_r [6] ? _12449_ : _12386_;
  assign _12451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [11] : \MSYNC_1r1w.synth.nz.mem[128] [11];
  assign _12452_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [11] : \MSYNC_1r1w.synth.nz.mem[130] [11];
  assign _12453_ = \bapg_rd.w_ptr_r [1] ? _12452_ : _12451_;
  assign _12454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [11] : \MSYNC_1r1w.synth.nz.mem[132] [11];
  assign _12455_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [11] : \MSYNC_1r1w.synth.nz.mem[134] [11];
  assign _12456_ = \bapg_rd.w_ptr_r [1] ? _12455_ : _12454_;
  assign _12457_ = \bapg_rd.w_ptr_r [2] ? _12456_ : _12453_;
  assign _12458_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [11] : \MSYNC_1r1w.synth.nz.mem[136] [11];
  assign _12459_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [11] : \MSYNC_1r1w.synth.nz.mem[138] [11];
  assign _12460_ = \bapg_rd.w_ptr_r [1] ? _12459_ : _12458_;
  assign _12461_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [11] : \MSYNC_1r1w.synth.nz.mem[140] [11];
  assign _12462_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [11] : \MSYNC_1r1w.synth.nz.mem[142] [11];
  assign _12463_ = \bapg_rd.w_ptr_r [1] ? _12462_ : _12461_;
  assign _12464_ = \bapg_rd.w_ptr_r [2] ? _12463_ : _12460_;
  assign _12465_ = \bapg_rd.w_ptr_r [3] ? _12464_ : _12457_;
  assign _12466_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [11] : \MSYNC_1r1w.synth.nz.mem[144] [11];
  assign _12467_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [11] : \MSYNC_1r1w.synth.nz.mem[146] [11];
  assign _12468_ = \bapg_rd.w_ptr_r [1] ? _12467_ : _12466_;
  assign _12469_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [11] : \MSYNC_1r1w.synth.nz.mem[148] [11];
  assign _12470_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [11] : \MSYNC_1r1w.synth.nz.mem[150] [11];
  assign _12471_ = \bapg_rd.w_ptr_r [1] ? _12470_ : _12469_;
  assign _12472_ = \bapg_rd.w_ptr_r [2] ? _12471_ : _12468_;
  assign _12473_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [11] : \MSYNC_1r1w.synth.nz.mem[152] [11];
  assign _12474_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [11] : \MSYNC_1r1w.synth.nz.mem[154] [11];
  assign _12475_ = \bapg_rd.w_ptr_r [1] ? _12474_ : _12473_;
  assign _12476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [11] : \MSYNC_1r1w.synth.nz.mem[156] [11];
  assign _12477_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [11] : \MSYNC_1r1w.synth.nz.mem[158] [11];
  assign _12478_ = \bapg_rd.w_ptr_r [1] ? _12477_ : _12476_;
  assign _12479_ = \bapg_rd.w_ptr_r [2] ? _12478_ : _12475_;
  assign _12480_ = \bapg_rd.w_ptr_r [3] ? _12479_ : _12472_;
  assign _12481_ = \bapg_rd.w_ptr_r [4] ? _12480_ : _12465_;
  assign _12482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [11] : \MSYNC_1r1w.synth.nz.mem[160] [11];
  assign _12483_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [11] : \MSYNC_1r1w.synth.nz.mem[162] [11];
  assign _12484_ = \bapg_rd.w_ptr_r [1] ? _12483_ : _12482_;
  assign _12485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [11] : \MSYNC_1r1w.synth.nz.mem[164] [11];
  assign _12486_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [11] : \MSYNC_1r1w.synth.nz.mem[166] [11];
  assign _12487_ = \bapg_rd.w_ptr_r [1] ? _12486_ : _12485_;
  assign _12488_ = \bapg_rd.w_ptr_r [2] ? _12487_ : _12484_;
  assign _12489_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [11] : \MSYNC_1r1w.synth.nz.mem[168] [11];
  assign _12490_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [11] : \MSYNC_1r1w.synth.nz.mem[170] [11];
  assign _12491_ = \bapg_rd.w_ptr_r [1] ? _12490_ : _12489_;
  assign _12492_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [11] : \MSYNC_1r1w.synth.nz.mem[172] [11];
  assign _12493_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [11] : \MSYNC_1r1w.synth.nz.mem[174] [11];
  assign _12494_ = \bapg_rd.w_ptr_r [1] ? _12493_ : _12492_;
  assign _12495_ = \bapg_rd.w_ptr_r [2] ? _12494_ : _12491_;
  assign _12496_ = \bapg_rd.w_ptr_r [3] ? _12495_ : _12488_;
  assign _12497_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [11] : \MSYNC_1r1w.synth.nz.mem[176] [11];
  assign _12498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [11] : \MSYNC_1r1w.synth.nz.mem[178] [11];
  assign _12499_ = \bapg_rd.w_ptr_r [1] ? _12498_ : _12497_;
  assign _12500_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [11] : \MSYNC_1r1w.synth.nz.mem[180] [11];
  assign _12501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [11] : \MSYNC_1r1w.synth.nz.mem[182] [11];
  assign _12502_ = \bapg_rd.w_ptr_r [1] ? _12501_ : _12500_;
  assign _12503_ = \bapg_rd.w_ptr_r [2] ? _12502_ : _12499_;
  assign _12504_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [11] : \MSYNC_1r1w.synth.nz.mem[184] [11];
  assign _12505_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [11] : \MSYNC_1r1w.synth.nz.mem[186] [11];
  assign _12506_ = \bapg_rd.w_ptr_r [1] ? _12505_ : _12504_;
  assign _12507_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [11] : \MSYNC_1r1w.synth.nz.mem[188] [11];
  assign _12508_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [11] : \MSYNC_1r1w.synth.nz.mem[190] [11];
  assign _12509_ = \bapg_rd.w_ptr_r [1] ? _12508_ : _12507_;
  assign _12510_ = \bapg_rd.w_ptr_r [2] ? _12509_ : _12506_;
  assign _12511_ = \bapg_rd.w_ptr_r [3] ? _12510_ : _12503_;
  assign _12512_ = \bapg_rd.w_ptr_r [4] ? _12511_ : _12496_;
  assign _12513_ = \bapg_rd.w_ptr_r [5] ? _12512_ : _12481_;
  assign _12514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [11] : \MSYNC_1r1w.synth.nz.mem[192] [11];
  assign _12515_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [11] : \MSYNC_1r1w.synth.nz.mem[194] [11];
  assign _12516_ = \bapg_rd.w_ptr_r [1] ? _12515_ : _12514_;
  assign _12517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [11] : \MSYNC_1r1w.synth.nz.mem[196] [11];
  assign _12518_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [11] : \MSYNC_1r1w.synth.nz.mem[198] [11];
  assign _12519_ = \bapg_rd.w_ptr_r [1] ? _12518_ : _12517_;
  assign _12520_ = \bapg_rd.w_ptr_r [2] ? _12519_ : _12516_;
  assign _12521_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [11] : \MSYNC_1r1w.synth.nz.mem[200] [11];
  assign _12522_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [11] : \MSYNC_1r1w.synth.nz.mem[202] [11];
  assign _12523_ = \bapg_rd.w_ptr_r [1] ? _12522_ : _12521_;
  assign _12524_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [11] : \MSYNC_1r1w.synth.nz.mem[204] [11];
  assign _12525_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [11] : \MSYNC_1r1w.synth.nz.mem[206] [11];
  assign _12526_ = \bapg_rd.w_ptr_r [1] ? _12525_ : _12524_;
  assign _12527_ = \bapg_rd.w_ptr_r [2] ? _12526_ : _12523_;
  assign _12528_ = \bapg_rd.w_ptr_r [3] ? _12527_ : _12520_;
  assign _12529_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [11] : \MSYNC_1r1w.synth.nz.mem[208] [11];
  assign _12530_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [11] : \MSYNC_1r1w.synth.nz.mem[210] [11];
  assign _12531_ = \bapg_rd.w_ptr_r [1] ? _12530_ : _12529_;
  assign _12532_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [11] : \MSYNC_1r1w.synth.nz.mem[212] [11];
  assign _12533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [11] : \MSYNC_1r1w.synth.nz.mem[214] [11];
  assign _12534_ = \bapg_rd.w_ptr_r [1] ? _12533_ : _12532_;
  assign _12535_ = \bapg_rd.w_ptr_r [2] ? _12534_ : _12531_;
  assign _12536_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [11] : \MSYNC_1r1w.synth.nz.mem[216] [11];
  assign _12537_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [11] : \MSYNC_1r1w.synth.nz.mem[218] [11];
  assign _12538_ = \bapg_rd.w_ptr_r [1] ? _12537_ : _12536_;
  assign _12539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [11] : \MSYNC_1r1w.synth.nz.mem[220] [11];
  assign _12540_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [11] : \MSYNC_1r1w.synth.nz.mem[222] [11];
  assign _12541_ = \bapg_rd.w_ptr_r [1] ? _12540_ : _12539_;
  assign _12542_ = \bapg_rd.w_ptr_r [2] ? _12541_ : _12538_;
  assign _12543_ = \bapg_rd.w_ptr_r [3] ? _12542_ : _12535_;
  assign _12544_ = \bapg_rd.w_ptr_r [4] ? _12543_ : _12528_;
  assign _12545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [11] : \MSYNC_1r1w.synth.nz.mem[224] [11];
  assign _12546_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [11] : \MSYNC_1r1w.synth.nz.mem[226] [11];
  assign _12547_ = \bapg_rd.w_ptr_r [1] ? _12546_ : _12545_;
  assign _12548_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [11] : \MSYNC_1r1w.synth.nz.mem[228] [11];
  assign _12549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [11] : \MSYNC_1r1w.synth.nz.mem[230] [11];
  assign _12550_ = \bapg_rd.w_ptr_r [1] ? _12549_ : _12548_;
  assign _12551_ = \bapg_rd.w_ptr_r [2] ? _12550_ : _12547_;
  assign _12552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [11] : \MSYNC_1r1w.synth.nz.mem[232] [11];
  assign _12553_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [11] : \MSYNC_1r1w.synth.nz.mem[234] [11];
  assign _12554_ = \bapg_rd.w_ptr_r [1] ? _12553_ : _12552_;
  assign _12555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [11] : \MSYNC_1r1w.synth.nz.mem[236] [11];
  assign _12556_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [11] : \MSYNC_1r1w.synth.nz.mem[238] [11];
  assign _12557_ = \bapg_rd.w_ptr_r [1] ? _12556_ : _12555_;
  assign _12558_ = \bapg_rd.w_ptr_r [2] ? _12557_ : _12554_;
  assign _12559_ = \bapg_rd.w_ptr_r [3] ? _12558_ : _12551_;
  assign _12560_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [11] : \MSYNC_1r1w.synth.nz.mem[240] [11];
  assign _12561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [11] : \MSYNC_1r1w.synth.nz.mem[242] [11];
  assign _12562_ = \bapg_rd.w_ptr_r [1] ? _12561_ : _12560_;
  assign _12563_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [11] : \MSYNC_1r1w.synth.nz.mem[244] [11];
  assign _12564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [11] : \MSYNC_1r1w.synth.nz.mem[246] [11];
  assign _12565_ = \bapg_rd.w_ptr_r [1] ? _12564_ : _12563_;
  assign _12566_ = \bapg_rd.w_ptr_r [2] ? _12565_ : _12562_;
  assign _12567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [11] : \MSYNC_1r1w.synth.nz.mem[248] [11];
  assign _12568_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [11] : \MSYNC_1r1w.synth.nz.mem[250] [11];
  assign _12569_ = \bapg_rd.w_ptr_r [1] ? _12568_ : _12567_;
  assign _12570_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [11] : \MSYNC_1r1w.synth.nz.mem[252] [11];
  assign _12571_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [11] : \MSYNC_1r1w.synth.nz.mem[254] [11];
  assign _12572_ = \bapg_rd.w_ptr_r [1] ? _12571_ : _12570_;
  assign _12573_ = \bapg_rd.w_ptr_r [2] ? _12572_ : _12569_;
  assign _12574_ = \bapg_rd.w_ptr_r [3] ? _12573_ : _12566_;
  assign _12575_ = \bapg_rd.w_ptr_r [4] ? _12574_ : _12559_;
  assign _12576_ = \bapg_rd.w_ptr_r [5] ? _12575_ : _12544_;
  assign _12577_ = \bapg_rd.w_ptr_r [6] ? _12576_ : _12513_;
  assign _12578_ = \bapg_rd.w_ptr_r [7] ? _12577_ : _12450_;
  assign _12579_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [11] : \MSYNC_1r1w.synth.nz.mem[256] [11];
  assign _12580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [11] : \MSYNC_1r1w.synth.nz.mem[258] [11];
  assign _12581_ = \bapg_rd.w_ptr_r [1] ? _12580_ : _12579_;
  assign _12582_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [11] : \MSYNC_1r1w.synth.nz.mem[260] [11];
  assign _12583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [11] : \MSYNC_1r1w.synth.nz.mem[262] [11];
  assign _12584_ = \bapg_rd.w_ptr_r [1] ? _12583_ : _12582_;
  assign _12585_ = \bapg_rd.w_ptr_r [2] ? _12584_ : _12581_;
  assign _12586_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [11] : \MSYNC_1r1w.synth.nz.mem[264] [11];
  assign _12587_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [11] : \MSYNC_1r1w.synth.nz.mem[266] [11];
  assign _12588_ = \bapg_rd.w_ptr_r [1] ? _12587_ : _12586_;
  assign _12589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [11] : \MSYNC_1r1w.synth.nz.mem[268] [11];
  assign _12590_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [11] : \MSYNC_1r1w.synth.nz.mem[270] [11];
  assign _12591_ = \bapg_rd.w_ptr_r [1] ? _12590_ : _12589_;
  assign _12592_ = \bapg_rd.w_ptr_r [2] ? _12591_ : _12588_;
  assign _12593_ = \bapg_rd.w_ptr_r [3] ? _12592_ : _12585_;
  assign _12594_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [11] : \MSYNC_1r1w.synth.nz.mem[272] [11];
  assign _12595_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [11] : \MSYNC_1r1w.synth.nz.mem[274] [11];
  assign _12596_ = \bapg_rd.w_ptr_r [1] ? _12595_ : _12594_;
  assign _12597_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [11] : \MSYNC_1r1w.synth.nz.mem[276] [11];
  assign _12598_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [11] : \MSYNC_1r1w.synth.nz.mem[278] [11];
  assign _12599_ = \bapg_rd.w_ptr_r [1] ? _12598_ : _12597_;
  assign _12600_ = \bapg_rd.w_ptr_r [2] ? _12599_ : _12596_;
  assign _12601_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [11] : \MSYNC_1r1w.synth.nz.mem[280] [11];
  assign _12602_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [11] : \MSYNC_1r1w.synth.nz.mem[282] [11];
  assign _12603_ = \bapg_rd.w_ptr_r [1] ? _12602_ : _12601_;
  assign _12604_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [11] : \MSYNC_1r1w.synth.nz.mem[284] [11];
  assign _12605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [11] : \MSYNC_1r1w.synth.nz.mem[286] [11];
  assign _12606_ = \bapg_rd.w_ptr_r [1] ? _12605_ : _12604_;
  assign _12607_ = \bapg_rd.w_ptr_r [2] ? _12606_ : _12603_;
  assign _12608_ = \bapg_rd.w_ptr_r [3] ? _12607_ : _12600_;
  assign _12609_ = \bapg_rd.w_ptr_r [4] ? _12608_ : _12593_;
  assign _12610_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [11] : \MSYNC_1r1w.synth.nz.mem[288] [11];
  assign _12611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [11] : \MSYNC_1r1w.synth.nz.mem[290] [11];
  assign _12612_ = \bapg_rd.w_ptr_r [1] ? _12611_ : _12610_;
  assign _12613_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [11] : \MSYNC_1r1w.synth.nz.mem[292] [11];
  assign _12614_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [11] : \MSYNC_1r1w.synth.nz.mem[294] [11];
  assign _12615_ = \bapg_rd.w_ptr_r [1] ? _12614_ : _12613_;
  assign _12616_ = \bapg_rd.w_ptr_r [2] ? _12615_ : _12612_;
  assign _12617_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [11] : \MSYNC_1r1w.synth.nz.mem[296] [11];
  assign _12618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [11] : \MSYNC_1r1w.synth.nz.mem[298] [11];
  assign _12619_ = \bapg_rd.w_ptr_r [1] ? _12618_ : _12617_;
  assign _12620_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [11] : \MSYNC_1r1w.synth.nz.mem[300] [11];
  assign _12621_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [11] : \MSYNC_1r1w.synth.nz.mem[302] [11];
  assign _12622_ = \bapg_rd.w_ptr_r [1] ? _12621_ : _12620_;
  assign _12623_ = \bapg_rd.w_ptr_r [2] ? _12622_ : _12619_;
  assign _12624_ = \bapg_rd.w_ptr_r [3] ? _12623_ : _12616_;
  assign _12625_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [11] : \MSYNC_1r1w.synth.nz.mem[304] [11];
  assign _12626_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [11] : \MSYNC_1r1w.synth.nz.mem[306] [11];
  assign _12627_ = \bapg_rd.w_ptr_r [1] ? _12626_ : _12625_;
  assign _12628_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [11] : \MSYNC_1r1w.synth.nz.mem[308] [11];
  assign _12629_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [11] : \MSYNC_1r1w.synth.nz.mem[310] [11];
  assign _12630_ = \bapg_rd.w_ptr_r [1] ? _12629_ : _12628_;
  assign _12631_ = \bapg_rd.w_ptr_r [2] ? _12630_ : _12627_;
  assign _12632_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [11] : \MSYNC_1r1w.synth.nz.mem[312] [11];
  assign _12633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [11] : \MSYNC_1r1w.synth.nz.mem[314] [11];
  assign _12634_ = \bapg_rd.w_ptr_r [1] ? _12633_ : _12632_;
  assign _12635_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [11] : \MSYNC_1r1w.synth.nz.mem[316] [11];
  assign _12636_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [11] : \MSYNC_1r1w.synth.nz.mem[318] [11];
  assign _12637_ = \bapg_rd.w_ptr_r [1] ? _12636_ : _12635_;
  assign _12638_ = \bapg_rd.w_ptr_r [2] ? _12637_ : _12634_;
  assign _12639_ = \bapg_rd.w_ptr_r [3] ? _12638_ : _12631_;
  assign _12640_ = \bapg_rd.w_ptr_r [4] ? _12639_ : _12624_;
  assign _12641_ = \bapg_rd.w_ptr_r [5] ? _12640_ : _12609_;
  assign _12642_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [11] : \MSYNC_1r1w.synth.nz.mem[320] [11];
  assign _12643_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [11] : \MSYNC_1r1w.synth.nz.mem[322] [11];
  assign _12644_ = \bapg_rd.w_ptr_r [1] ? _12643_ : _12642_;
  assign _12645_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [11] : \MSYNC_1r1w.synth.nz.mem[324] [11];
  assign _12646_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [11] : \MSYNC_1r1w.synth.nz.mem[326] [11];
  assign _12647_ = \bapg_rd.w_ptr_r [1] ? _12646_ : _12645_;
  assign _12648_ = \bapg_rd.w_ptr_r [2] ? _12647_ : _12644_;
  assign _12649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [11] : \MSYNC_1r1w.synth.nz.mem[328] [11];
  assign _12650_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [11] : \MSYNC_1r1w.synth.nz.mem[330] [11];
  assign _12651_ = \bapg_rd.w_ptr_r [1] ? _12650_ : _12649_;
  assign _12652_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [11] : \MSYNC_1r1w.synth.nz.mem[332] [11];
  assign _12653_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [11] : \MSYNC_1r1w.synth.nz.mem[334] [11];
  assign _12654_ = \bapg_rd.w_ptr_r [1] ? _12653_ : _12652_;
  assign _12655_ = \bapg_rd.w_ptr_r [2] ? _12654_ : _12651_;
  assign _12656_ = \bapg_rd.w_ptr_r [3] ? _12655_ : _12648_;
  assign _12657_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [11] : \MSYNC_1r1w.synth.nz.mem[336] [11];
  assign _12658_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [11] : \MSYNC_1r1w.synth.nz.mem[338] [11];
  assign _12659_ = \bapg_rd.w_ptr_r [1] ? _12658_ : _12657_;
  assign _12660_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [11] : \MSYNC_1r1w.synth.nz.mem[340] [11];
  assign _12661_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [11] : \MSYNC_1r1w.synth.nz.mem[342] [11];
  assign _12662_ = \bapg_rd.w_ptr_r [1] ? _12661_ : _12660_;
  assign _12663_ = \bapg_rd.w_ptr_r [2] ? _12662_ : _12659_;
  assign _12664_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [11] : \MSYNC_1r1w.synth.nz.mem[344] [11];
  assign _12665_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [11] : \MSYNC_1r1w.synth.nz.mem[346] [11];
  assign _12666_ = \bapg_rd.w_ptr_r [1] ? _12665_ : _12664_;
  assign _12667_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [11] : \MSYNC_1r1w.synth.nz.mem[348] [11];
  assign _12668_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [11] : \MSYNC_1r1w.synth.nz.mem[350] [11];
  assign _12669_ = \bapg_rd.w_ptr_r [1] ? _12668_ : _12667_;
  assign _12670_ = \bapg_rd.w_ptr_r [2] ? _12669_ : _12666_;
  assign _12671_ = \bapg_rd.w_ptr_r [3] ? _12670_ : _12663_;
  assign _12672_ = \bapg_rd.w_ptr_r [4] ? _12671_ : _12656_;
  assign _12673_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [11] : \MSYNC_1r1w.synth.nz.mem[352] [11];
  assign _12674_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [11] : \MSYNC_1r1w.synth.nz.mem[354] [11];
  assign _12675_ = \bapg_rd.w_ptr_r [1] ? _12674_ : _12673_;
  assign _12676_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [11] : \MSYNC_1r1w.synth.nz.mem[356] [11];
  assign _12677_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [11] : \MSYNC_1r1w.synth.nz.mem[358] [11];
  assign _12678_ = \bapg_rd.w_ptr_r [1] ? _12677_ : _12676_;
  assign _12679_ = \bapg_rd.w_ptr_r [2] ? _12678_ : _12675_;
  assign _12680_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [11] : \MSYNC_1r1w.synth.nz.mem[360] [11];
  assign _12681_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [11] : \MSYNC_1r1w.synth.nz.mem[362] [11];
  assign _12682_ = \bapg_rd.w_ptr_r [1] ? _12681_ : _12680_;
  assign _12683_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [11] : \MSYNC_1r1w.synth.nz.mem[364] [11];
  assign _12684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [11] : \MSYNC_1r1w.synth.nz.mem[366] [11];
  assign _12685_ = \bapg_rd.w_ptr_r [1] ? _12684_ : _12683_;
  assign _12686_ = \bapg_rd.w_ptr_r [2] ? _12685_ : _12682_;
  assign _12687_ = \bapg_rd.w_ptr_r [3] ? _12686_ : _12679_;
  assign _12688_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [11] : \MSYNC_1r1w.synth.nz.mem[368] [11];
  assign _12689_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [11] : \MSYNC_1r1w.synth.nz.mem[370] [11];
  assign _12690_ = \bapg_rd.w_ptr_r [1] ? _12689_ : _12688_;
  assign _12691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [11] : \MSYNC_1r1w.synth.nz.mem[372] [11];
  assign _12692_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [11] : \MSYNC_1r1w.synth.nz.mem[374] [11];
  assign _12693_ = \bapg_rd.w_ptr_r [1] ? _12692_ : _12691_;
  assign _12694_ = \bapg_rd.w_ptr_r [2] ? _12693_ : _12690_;
  assign _12695_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [11] : \MSYNC_1r1w.synth.nz.mem[376] [11];
  assign _12696_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [11] : \MSYNC_1r1w.synth.nz.mem[378] [11];
  assign _12697_ = \bapg_rd.w_ptr_r [1] ? _12696_ : _12695_;
  assign _12698_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [11] : \MSYNC_1r1w.synth.nz.mem[380] [11];
  assign _12699_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [11] : \MSYNC_1r1w.synth.nz.mem[382] [11];
  assign _12700_ = \bapg_rd.w_ptr_r [1] ? _12699_ : _12698_;
  assign _12701_ = \bapg_rd.w_ptr_r [2] ? _12700_ : _12697_;
  assign _12702_ = \bapg_rd.w_ptr_r [3] ? _12701_ : _12694_;
  assign _12703_ = \bapg_rd.w_ptr_r [4] ? _12702_ : _12687_;
  assign _12704_ = \bapg_rd.w_ptr_r [5] ? _12703_ : _12672_;
  assign _12705_ = \bapg_rd.w_ptr_r [6] ? _12704_ : _12641_;
  assign _12706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [11] : \MSYNC_1r1w.synth.nz.mem[384] [11];
  assign _12707_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [11] : \MSYNC_1r1w.synth.nz.mem[386] [11];
  assign _12708_ = \bapg_rd.w_ptr_r [1] ? _12707_ : _12706_;
  assign _12709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [11] : \MSYNC_1r1w.synth.nz.mem[388] [11];
  assign _12710_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [11] : \MSYNC_1r1w.synth.nz.mem[390] [11];
  assign _12711_ = \bapg_rd.w_ptr_r [1] ? _12710_ : _12709_;
  assign _12712_ = \bapg_rd.w_ptr_r [2] ? _12711_ : _12708_;
  assign _12713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [11] : \MSYNC_1r1w.synth.nz.mem[392] [11];
  assign _12714_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [11] : \MSYNC_1r1w.synth.nz.mem[394] [11];
  assign _12715_ = \bapg_rd.w_ptr_r [1] ? _12714_ : _12713_;
  assign _12716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [11] : \MSYNC_1r1w.synth.nz.mem[396] [11];
  assign _12717_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [11] : \MSYNC_1r1w.synth.nz.mem[398] [11];
  assign _12718_ = \bapg_rd.w_ptr_r [1] ? _12717_ : _12716_;
  assign _12719_ = \bapg_rd.w_ptr_r [2] ? _12718_ : _12715_;
  assign _12720_ = \bapg_rd.w_ptr_r [3] ? _12719_ : _12712_;
  assign _12721_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [11] : \MSYNC_1r1w.synth.nz.mem[400] [11];
  assign _12722_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [11] : \MSYNC_1r1w.synth.nz.mem[402] [11];
  assign _12723_ = \bapg_rd.w_ptr_r [1] ? _12722_ : _12721_;
  assign _12724_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [11] : \MSYNC_1r1w.synth.nz.mem[404] [11];
  assign _12725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [11] : \MSYNC_1r1w.synth.nz.mem[406] [11];
  assign _12726_ = \bapg_rd.w_ptr_r [1] ? _12725_ : _12724_;
  assign _12727_ = \bapg_rd.w_ptr_r [2] ? _12726_ : _12723_;
  assign _12728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [11] : \MSYNC_1r1w.synth.nz.mem[408] [11];
  assign _12729_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [11] : \MSYNC_1r1w.synth.nz.mem[410] [11];
  assign _12730_ = \bapg_rd.w_ptr_r [1] ? _12729_ : _12728_;
  assign _12731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [11] : \MSYNC_1r1w.synth.nz.mem[412] [11];
  assign _12732_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [11] : \MSYNC_1r1w.synth.nz.mem[414] [11];
  assign _12733_ = \bapg_rd.w_ptr_r [1] ? _12732_ : _12731_;
  assign _12734_ = \bapg_rd.w_ptr_r [2] ? _12733_ : _12730_;
  assign _12735_ = \bapg_rd.w_ptr_r [3] ? _12734_ : _12727_;
  assign _12736_ = \bapg_rd.w_ptr_r [4] ? _12735_ : _12720_;
  assign _12737_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [11] : \MSYNC_1r1w.synth.nz.mem[416] [11];
  assign _12738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [11] : \MSYNC_1r1w.synth.nz.mem[418] [11];
  assign _12739_ = \bapg_rd.w_ptr_r [1] ? _12738_ : _12737_;
  assign _12740_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [11] : \MSYNC_1r1w.synth.nz.mem[420] [11];
  assign _12741_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [11] : \MSYNC_1r1w.synth.nz.mem[422] [11];
  assign _12742_ = \bapg_rd.w_ptr_r [1] ? _12741_ : _12740_;
  assign _12743_ = \bapg_rd.w_ptr_r [2] ? _12742_ : _12739_;
  assign _12744_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [11] : \MSYNC_1r1w.synth.nz.mem[424] [11];
  assign _12745_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [11] : \MSYNC_1r1w.synth.nz.mem[426] [11];
  assign _12746_ = \bapg_rd.w_ptr_r [1] ? _12745_ : _12744_;
  assign _12747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [11] : \MSYNC_1r1w.synth.nz.mem[428] [11];
  assign _12748_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [11] : \MSYNC_1r1w.synth.nz.mem[430] [11];
  assign _12749_ = \bapg_rd.w_ptr_r [1] ? _12748_ : _12747_;
  assign _12750_ = \bapg_rd.w_ptr_r [2] ? _12749_ : _12746_;
  assign _12751_ = \bapg_rd.w_ptr_r [3] ? _12750_ : _12743_;
  assign _12752_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [11] : \MSYNC_1r1w.synth.nz.mem[432] [11];
  assign _12753_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [11] : \MSYNC_1r1w.synth.nz.mem[434] [11];
  assign _12754_ = \bapg_rd.w_ptr_r [1] ? _12753_ : _12752_;
  assign _12755_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [11] : \MSYNC_1r1w.synth.nz.mem[436] [11];
  assign _12756_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [11] : \MSYNC_1r1w.synth.nz.mem[438] [11];
  assign _12757_ = \bapg_rd.w_ptr_r [1] ? _12756_ : _12755_;
  assign _12758_ = \bapg_rd.w_ptr_r [2] ? _12757_ : _12754_;
  assign _12759_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [11] : \MSYNC_1r1w.synth.nz.mem[440] [11];
  assign _12760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [11] : \MSYNC_1r1w.synth.nz.mem[442] [11];
  assign _12761_ = \bapg_rd.w_ptr_r [1] ? _12760_ : _12759_;
  assign _12762_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [11] : \MSYNC_1r1w.synth.nz.mem[444] [11];
  assign _12763_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [11] : \MSYNC_1r1w.synth.nz.mem[446] [11];
  assign _12764_ = \bapg_rd.w_ptr_r [1] ? _12763_ : _12762_;
  assign _12765_ = \bapg_rd.w_ptr_r [2] ? _12764_ : _12761_;
  assign _12766_ = \bapg_rd.w_ptr_r [3] ? _12765_ : _12758_;
  assign _12767_ = \bapg_rd.w_ptr_r [4] ? _12766_ : _12751_;
  assign _12768_ = \bapg_rd.w_ptr_r [5] ? _12767_ : _12736_;
  assign _12769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [11] : \MSYNC_1r1w.synth.nz.mem[448] [11];
  assign _12770_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [11] : \MSYNC_1r1w.synth.nz.mem[450] [11];
  assign _12771_ = \bapg_rd.w_ptr_r [1] ? _12770_ : _12769_;
  assign _12772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [11] : \MSYNC_1r1w.synth.nz.mem[452] [11];
  assign _12773_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [11] : \MSYNC_1r1w.synth.nz.mem[454] [11];
  assign _12774_ = \bapg_rd.w_ptr_r [1] ? _12773_ : _12772_;
  assign _12775_ = \bapg_rd.w_ptr_r [2] ? _12774_ : _12771_;
  assign _12776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [11] : \MSYNC_1r1w.synth.nz.mem[456] [11];
  assign _12777_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [11] : \MSYNC_1r1w.synth.nz.mem[458] [11];
  assign _12778_ = \bapg_rd.w_ptr_r [1] ? _12777_ : _12776_;
  assign _12779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [11] : \MSYNC_1r1w.synth.nz.mem[460] [11];
  assign _12780_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [11] : \MSYNC_1r1w.synth.nz.mem[462] [11];
  assign _12781_ = \bapg_rd.w_ptr_r [1] ? _12780_ : _12779_;
  assign _12782_ = \bapg_rd.w_ptr_r [2] ? _12781_ : _12778_;
  assign _12783_ = \bapg_rd.w_ptr_r [3] ? _12782_ : _12775_;
  assign _12784_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [11] : \MSYNC_1r1w.synth.nz.mem[464] [11];
  assign _12785_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [11] : \MSYNC_1r1w.synth.nz.mem[466] [11];
  assign _12786_ = \bapg_rd.w_ptr_r [1] ? _12785_ : _12784_;
  assign _12787_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [11] : \MSYNC_1r1w.synth.nz.mem[468] [11];
  assign _12788_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [11] : \MSYNC_1r1w.synth.nz.mem[470] [11];
  assign _12789_ = \bapg_rd.w_ptr_r [1] ? _12788_ : _12787_;
  assign _12790_ = \bapg_rd.w_ptr_r [2] ? _12789_ : _12786_;
  assign _12791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [11] : \MSYNC_1r1w.synth.nz.mem[472] [11];
  assign _12792_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [11] : \MSYNC_1r1w.synth.nz.mem[474] [11];
  assign _12793_ = \bapg_rd.w_ptr_r [1] ? _12792_ : _12791_;
  assign _12794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [11] : \MSYNC_1r1w.synth.nz.mem[476] [11];
  assign _12795_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [11] : \MSYNC_1r1w.synth.nz.mem[478] [11];
  assign _12796_ = \bapg_rd.w_ptr_r [1] ? _12795_ : _12794_;
  assign _12797_ = \bapg_rd.w_ptr_r [2] ? _12796_ : _12793_;
  assign _12798_ = \bapg_rd.w_ptr_r [3] ? _12797_ : _12790_;
  assign _12799_ = \bapg_rd.w_ptr_r [4] ? _12798_ : _12783_;
  assign _12800_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [11] : \MSYNC_1r1w.synth.nz.mem[480] [11];
  assign _12801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [11] : \MSYNC_1r1w.synth.nz.mem[482] [11];
  assign _12802_ = \bapg_rd.w_ptr_r [1] ? _12801_ : _12800_;
  assign _12803_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [11] : \MSYNC_1r1w.synth.nz.mem[484] [11];
  assign _12804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [11] : \MSYNC_1r1w.synth.nz.mem[486] [11];
  assign _12805_ = \bapg_rd.w_ptr_r [1] ? _12804_ : _12803_;
  assign _12806_ = \bapg_rd.w_ptr_r [2] ? _12805_ : _12802_;
  assign _12807_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [11] : \MSYNC_1r1w.synth.nz.mem[488] [11];
  assign _12808_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [11] : \MSYNC_1r1w.synth.nz.mem[490] [11];
  assign _12809_ = \bapg_rd.w_ptr_r [1] ? _12808_ : _12807_;
  assign _12810_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [11] : \MSYNC_1r1w.synth.nz.mem[492] [11];
  assign _12811_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [11] : \MSYNC_1r1w.synth.nz.mem[494] [11];
  assign _12812_ = \bapg_rd.w_ptr_r [1] ? _12811_ : _12810_;
  assign _12813_ = \bapg_rd.w_ptr_r [2] ? _12812_ : _12809_;
  assign _12814_ = \bapg_rd.w_ptr_r [3] ? _12813_ : _12806_;
  assign _12815_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [11] : \MSYNC_1r1w.synth.nz.mem[496] [11];
  assign _12816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [11] : \MSYNC_1r1w.synth.nz.mem[498] [11];
  assign _12817_ = \bapg_rd.w_ptr_r [1] ? _12816_ : _12815_;
  assign _12818_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [11] : \MSYNC_1r1w.synth.nz.mem[500] [11];
  assign _12819_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [11] : \MSYNC_1r1w.synth.nz.mem[502] [11];
  assign _12820_ = \bapg_rd.w_ptr_r [1] ? _12819_ : _12818_;
  assign _12821_ = \bapg_rd.w_ptr_r [2] ? _12820_ : _12817_;
  assign _12822_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [11] : \MSYNC_1r1w.synth.nz.mem[504] [11];
  assign _12823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [11] : \MSYNC_1r1w.synth.nz.mem[506] [11];
  assign _12824_ = \bapg_rd.w_ptr_r [1] ? _12823_ : _12822_;
  assign _12825_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [11] : \MSYNC_1r1w.synth.nz.mem[508] [11];
  assign _12826_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [11] : \MSYNC_1r1w.synth.nz.mem[510] [11];
  assign _12827_ = \bapg_rd.w_ptr_r [1] ? _12826_ : _12825_;
  assign _12828_ = \bapg_rd.w_ptr_r [2] ? _12827_ : _12824_;
  assign _12829_ = \bapg_rd.w_ptr_r [3] ? _12828_ : _12821_;
  assign _12830_ = \bapg_rd.w_ptr_r [4] ? _12829_ : _12814_;
  assign _12831_ = \bapg_rd.w_ptr_r [5] ? _12830_ : _12799_;
  assign _12832_ = \bapg_rd.w_ptr_r [6] ? _12831_ : _12768_;
  assign _12833_ = \bapg_rd.w_ptr_r [7] ? _12832_ : _12705_;
  assign _12834_ = \bapg_rd.w_ptr_r [8] ? _12833_ : _12578_;
  assign _12835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [11] : \MSYNC_1r1w.synth.nz.mem[512] [11];
  assign _12836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [11] : \MSYNC_1r1w.synth.nz.mem[514] [11];
  assign _12837_ = \bapg_rd.w_ptr_r [1] ? _12836_ : _12835_;
  assign _12838_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [11] : \MSYNC_1r1w.synth.nz.mem[516] [11];
  assign _12839_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [11] : \MSYNC_1r1w.synth.nz.mem[518] [11];
  assign _12840_ = \bapg_rd.w_ptr_r [1] ? _12839_ : _12838_;
  assign _12841_ = \bapg_rd.w_ptr_r [2] ? _12840_ : _12837_;
  assign _12842_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [11] : \MSYNC_1r1w.synth.nz.mem[520] [11];
  assign _12843_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [11] : \MSYNC_1r1w.synth.nz.mem[522] [11];
  assign _12844_ = \bapg_rd.w_ptr_r [1] ? _12843_ : _12842_;
  assign _12845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [11] : \MSYNC_1r1w.synth.nz.mem[524] [11];
  assign _12846_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [11] : \MSYNC_1r1w.synth.nz.mem[526] [11];
  assign _12847_ = \bapg_rd.w_ptr_r [1] ? _12846_ : _12845_;
  assign _12848_ = \bapg_rd.w_ptr_r [2] ? _12847_ : _12844_;
  assign _12849_ = \bapg_rd.w_ptr_r [3] ? _12848_ : _12841_;
  assign _12850_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [11] : \MSYNC_1r1w.synth.nz.mem[528] [11];
  assign _12851_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [11] : \MSYNC_1r1w.synth.nz.mem[530] [11];
  assign _12852_ = \bapg_rd.w_ptr_r [1] ? _12851_ : _12850_;
  assign _12853_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [11] : \MSYNC_1r1w.synth.nz.mem[532] [11];
  assign _12854_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [11] : \MSYNC_1r1w.synth.nz.mem[534] [11];
  assign _12855_ = \bapg_rd.w_ptr_r [1] ? _12854_ : _12853_;
  assign _12856_ = \bapg_rd.w_ptr_r [2] ? _12855_ : _12852_;
  assign _12857_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [11] : \MSYNC_1r1w.synth.nz.mem[536] [11];
  assign _12858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [11] : \MSYNC_1r1w.synth.nz.mem[538] [11];
  assign _12859_ = \bapg_rd.w_ptr_r [1] ? _12858_ : _12857_;
  assign _12860_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [11] : \MSYNC_1r1w.synth.nz.mem[540] [11];
  assign _12861_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [11] : \MSYNC_1r1w.synth.nz.mem[542] [11];
  assign _12862_ = \bapg_rd.w_ptr_r [1] ? _12861_ : _12860_;
  assign _12863_ = \bapg_rd.w_ptr_r [2] ? _12862_ : _12859_;
  assign _12864_ = \bapg_rd.w_ptr_r [3] ? _12863_ : _12856_;
  assign _12865_ = \bapg_rd.w_ptr_r [4] ? _12864_ : _12849_;
  assign _12866_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [11] : \MSYNC_1r1w.synth.nz.mem[544] [11];
  assign _12867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [11] : \MSYNC_1r1w.synth.nz.mem[546] [11];
  assign _12868_ = \bapg_rd.w_ptr_r [1] ? _12867_ : _12866_;
  assign _12869_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [11] : \MSYNC_1r1w.synth.nz.mem[548] [11];
  assign _12870_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [11] : \MSYNC_1r1w.synth.nz.mem[550] [11];
  assign _12871_ = \bapg_rd.w_ptr_r [1] ? _12870_ : _12869_;
  assign _12872_ = \bapg_rd.w_ptr_r [2] ? _12871_ : _12868_;
  assign _12873_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [11] : \MSYNC_1r1w.synth.nz.mem[552] [11];
  assign _12874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [11] : \MSYNC_1r1w.synth.nz.mem[554] [11];
  assign _12875_ = \bapg_rd.w_ptr_r [1] ? _12874_ : _12873_;
  assign _12876_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [11] : \MSYNC_1r1w.synth.nz.mem[556] [11];
  assign _12877_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [11] : \MSYNC_1r1w.synth.nz.mem[558] [11];
  assign _12878_ = \bapg_rd.w_ptr_r [1] ? _12877_ : _12876_;
  assign _12879_ = \bapg_rd.w_ptr_r [2] ? _12878_ : _12875_;
  assign _12880_ = \bapg_rd.w_ptr_r [3] ? _12879_ : _12872_;
  assign _12881_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [11] : \MSYNC_1r1w.synth.nz.mem[560] [11];
  assign _12882_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [11] : \MSYNC_1r1w.synth.nz.mem[562] [11];
  assign _12883_ = \bapg_rd.w_ptr_r [1] ? _12882_ : _12881_;
  assign _12884_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [11] : \MSYNC_1r1w.synth.nz.mem[564] [11];
  assign _12885_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [11] : \MSYNC_1r1w.synth.nz.mem[566] [11];
  assign _12886_ = \bapg_rd.w_ptr_r [1] ? _12885_ : _12884_;
  assign _12887_ = \bapg_rd.w_ptr_r [2] ? _12886_ : _12883_;
  assign _12888_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [11] : \MSYNC_1r1w.synth.nz.mem[568] [11];
  assign _12889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [11] : \MSYNC_1r1w.synth.nz.mem[570] [11];
  assign _12890_ = \bapg_rd.w_ptr_r [1] ? _12889_ : _12888_;
  assign _12891_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [11] : \MSYNC_1r1w.synth.nz.mem[572] [11];
  assign _12892_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [11] : \MSYNC_1r1w.synth.nz.mem[574] [11];
  assign _12893_ = \bapg_rd.w_ptr_r [1] ? _12892_ : _12891_;
  assign _12894_ = \bapg_rd.w_ptr_r [2] ? _12893_ : _12890_;
  assign _12895_ = \bapg_rd.w_ptr_r [3] ? _12894_ : _12887_;
  assign _12896_ = \bapg_rd.w_ptr_r [4] ? _12895_ : _12880_;
  assign _12897_ = \bapg_rd.w_ptr_r [5] ? _12896_ : _12865_;
  assign _12898_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [11] : \MSYNC_1r1w.synth.nz.mem[576] [11];
  assign _12899_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [11] : \MSYNC_1r1w.synth.nz.mem[578] [11];
  assign _12900_ = \bapg_rd.w_ptr_r [1] ? _12899_ : _12898_;
  assign _12901_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [11] : \MSYNC_1r1w.synth.nz.mem[580] [11];
  assign _12902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [11] : \MSYNC_1r1w.synth.nz.mem[582] [11];
  assign _12903_ = \bapg_rd.w_ptr_r [1] ? _12902_ : _12901_;
  assign _12904_ = \bapg_rd.w_ptr_r [2] ? _12903_ : _12900_;
  assign _12905_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [11] : \MSYNC_1r1w.synth.nz.mem[584] [11];
  assign _12906_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [11] : \MSYNC_1r1w.synth.nz.mem[586] [11];
  assign _12907_ = \bapg_rd.w_ptr_r [1] ? _12906_ : _12905_;
  assign _12908_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [11] : \MSYNC_1r1w.synth.nz.mem[588] [11];
  assign _12909_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [11] : \MSYNC_1r1w.synth.nz.mem[590] [11];
  assign _12910_ = \bapg_rd.w_ptr_r [1] ? _12909_ : _12908_;
  assign _12911_ = \bapg_rd.w_ptr_r [2] ? _12910_ : _12907_;
  assign _12912_ = \bapg_rd.w_ptr_r [3] ? _12911_ : _12904_;
  assign _12913_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [11] : \MSYNC_1r1w.synth.nz.mem[592] [11];
  assign _12914_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [11] : \MSYNC_1r1w.synth.nz.mem[594] [11];
  assign _12915_ = \bapg_rd.w_ptr_r [1] ? _12914_ : _12913_;
  assign _12916_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [11] : \MSYNC_1r1w.synth.nz.mem[596] [11];
  assign _12917_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [11] : \MSYNC_1r1w.synth.nz.mem[598] [11];
  assign _12918_ = \bapg_rd.w_ptr_r [1] ? _12917_ : _12916_;
  assign _12919_ = \bapg_rd.w_ptr_r [2] ? _12918_ : _12915_;
  assign _12920_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [11] : \MSYNC_1r1w.synth.nz.mem[600] [11];
  assign _12921_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [11] : \MSYNC_1r1w.synth.nz.mem[602] [11];
  assign _12922_ = \bapg_rd.w_ptr_r [1] ? _12921_ : _12920_;
  assign _12923_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [11] : \MSYNC_1r1w.synth.nz.mem[604] [11];
  assign _12924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [11] : \MSYNC_1r1w.synth.nz.mem[606] [11];
  assign _12925_ = \bapg_rd.w_ptr_r [1] ? _12924_ : _12923_;
  assign _12926_ = \bapg_rd.w_ptr_r [2] ? _12925_ : _12922_;
  assign _12927_ = \bapg_rd.w_ptr_r [3] ? _12926_ : _12919_;
  assign _12928_ = \bapg_rd.w_ptr_r [4] ? _12927_ : _12912_;
  assign _12929_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [11] : \MSYNC_1r1w.synth.nz.mem[608] [11];
  assign _12930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [11] : \MSYNC_1r1w.synth.nz.mem[610] [11];
  assign _12931_ = \bapg_rd.w_ptr_r [1] ? _12930_ : _12929_;
  assign _12932_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [11] : \MSYNC_1r1w.synth.nz.mem[612] [11];
  assign _12933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [11] : \MSYNC_1r1w.synth.nz.mem[614] [11];
  assign _12934_ = \bapg_rd.w_ptr_r [1] ? _12933_ : _12932_;
  assign _12935_ = \bapg_rd.w_ptr_r [2] ? _12934_ : _12931_;
  assign _12936_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [11] : \MSYNC_1r1w.synth.nz.mem[616] [11];
  assign _12937_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [11] : \MSYNC_1r1w.synth.nz.mem[618] [11];
  assign _12938_ = \bapg_rd.w_ptr_r [1] ? _12937_ : _12936_;
  assign _12939_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [11] : \MSYNC_1r1w.synth.nz.mem[620] [11];
  assign _12940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [11] : \MSYNC_1r1w.synth.nz.mem[622] [11];
  assign _12941_ = \bapg_rd.w_ptr_r [1] ? _12940_ : _12939_;
  assign _12942_ = \bapg_rd.w_ptr_r [2] ? _12941_ : _12938_;
  assign _12943_ = \bapg_rd.w_ptr_r [3] ? _12942_ : _12935_;
  assign _12944_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [11] : \MSYNC_1r1w.synth.nz.mem[624] [11];
  assign _12945_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [11] : \MSYNC_1r1w.synth.nz.mem[626] [11];
  assign _12946_ = \bapg_rd.w_ptr_r [1] ? _12945_ : _12944_;
  assign _12947_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [11] : \MSYNC_1r1w.synth.nz.mem[628] [11];
  assign _12948_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [11] : \MSYNC_1r1w.synth.nz.mem[630] [11];
  assign _12949_ = \bapg_rd.w_ptr_r [1] ? _12948_ : _12947_;
  assign _12950_ = \bapg_rd.w_ptr_r [2] ? _12949_ : _12946_;
  assign _12951_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [11] : \MSYNC_1r1w.synth.nz.mem[632] [11];
  assign _12952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [11] : \MSYNC_1r1w.synth.nz.mem[634] [11];
  assign _12953_ = \bapg_rd.w_ptr_r [1] ? _12952_ : _12951_;
  assign _12954_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [11] : \MSYNC_1r1w.synth.nz.mem[636] [11];
  assign _12955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [11] : \MSYNC_1r1w.synth.nz.mem[638] [11];
  assign _12956_ = \bapg_rd.w_ptr_r [1] ? _12955_ : _12954_;
  assign _12957_ = \bapg_rd.w_ptr_r [2] ? _12956_ : _12953_;
  assign _12958_ = \bapg_rd.w_ptr_r [3] ? _12957_ : _12950_;
  assign _12959_ = \bapg_rd.w_ptr_r [4] ? _12958_ : _12943_;
  assign _12960_ = \bapg_rd.w_ptr_r [5] ? _12959_ : _12928_;
  assign _12961_ = \bapg_rd.w_ptr_r [6] ? _12960_ : _12897_;
  assign _12962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [11] : \MSYNC_1r1w.synth.nz.mem[640] [11];
  assign _12963_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [11] : \MSYNC_1r1w.synth.nz.mem[642] [11];
  assign _12964_ = \bapg_rd.w_ptr_r [1] ? _12963_ : _12962_;
  assign _12965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [11] : \MSYNC_1r1w.synth.nz.mem[644] [11];
  assign _12966_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [11] : \MSYNC_1r1w.synth.nz.mem[646] [11];
  assign _12967_ = \bapg_rd.w_ptr_r [1] ? _12966_ : _12965_;
  assign _12968_ = \bapg_rd.w_ptr_r [2] ? _12967_ : _12964_;
  assign _12969_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [11] : \MSYNC_1r1w.synth.nz.mem[648] [11];
  assign _12970_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [11] : \MSYNC_1r1w.synth.nz.mem[650] [11];
  assign _12971_ = \bapg_rd.w_ptr_r [1] ? _12970_ : _12969_;
  assign _12972_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [11] : \MSYNC_1r1w.synth.nz.mem[652] [11];
  assign _12973_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [11] : \MSYNC_1r1w.synth.nz.mem[654] [11];
  assign _12974_ = \bapg_rd.w_ptr_r [1] ? _12973_ : _12972_;
  assign _12975_ = \bapg_rd.w_ptr_r [2] ? _12974_ : _12971_;
  assign _12976_ = \bapg_rd.w_ptr_r [3] ? _12975_ : _12968_;
  assign _12977_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [11] : \MSYNC_1r1w.synth.nz.mem[656] [11];
  assign _12978_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [11] : \MSYNC_1r1w.synth.nz.mem[658] [11];
  assign _12979_ = \bapg_rd.w_ptr_r [1] ? _12978_ : _12977_;
  assign _12980_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [11] : \MSYNC_1r1w.synth.nz.mem[660] [11];
  assign _12981_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [11] : \MSYNC_1r1w.synth.nz.mem[662] [11];
  assign _12982_ = \bapg_rd.w_ptr_r [1] ? _12981_ : _12980_;
  assign _12983_ = \bapg_rd.w_ptr_r [2] ? _12982_ : _12979_;
  assign _12984_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [11] : \MSYNC_1r1w.synth.nz.mem[664] [11];
  assign _12985_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [11] : \MSYNC_1r1w.synth.nz.mem[666] [11];
  assign _12986_ = \bapg_rd.w_ptr_r [1] ? _12985_ : _12984_;
  assign _12987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [11] : \MSYNC_1r1w.synth.nz.mem[668] [11];
  assign _12988_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [11] : \MSYNC_1r1w.synth.nz.mem[670] [11];
  assign _12989_ = \bapg_rd.w_ptr_r [1] ? _12988_ : _12987_;
  assign _12990_ = \bapg_rd.w_ptr_r [2] ? _12989_ : _12986_;
  assign _12991_ = \bapg_rd.w_ptr_r [3] ? _12990_ : _12983_;
  assign _12992_ = \bapg_rd.w_ptr_r [4] ? _12991_ : _12976_;
  assign _12993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [11] : \MSYNC_1r1w.synth.nz.mem[672] [11];
  assign _12994_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [11] : \MSYNC_1r1w.synth.nz.mem[674] [11];
  assign _12995_ = \bapg_rd.w_ptr_r [1] ? _12994_ : _12993_;
  assign _12996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [11] : \MSYNC_1r1w.synth.nz.mem[676] [11];
  assign _12997_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [11] : \MSYNC_1r1w.synth.nz.mem[678] [11];
  assign _12998_ = \bapg_rd.w_ptr_r [1] ? _12997_ : _12996_;
  assign _12999_ = \bapg_rd.w_ptr_r [2] ? _12998_ : _12995_;
  assign _13000_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [11] : \MSYNC_1r1w.synth.nz.mem[680] [11];
  assign _13001_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [11] : \MSYNC_1r1w.synth.nz.mem[682] [11];
  assign _13002_ = \bapg_rd.w_ptr_r [1] ? _13001_ : _13000_;
  assign _13003_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [11] : \MSYNC_1r1w.synth.nz.mem[684] [11];
  assign _13004_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [11] : \MSYNC_1r1w.synth.nz.mem[686] [11];
  assign _13005_ = \bapg_rd.w_ptr_r [1] ? _13004_ : _13003_;
  assign _13006_ = \bapg_rd.w_ptr_r [2] ? _13005_ : _13002_;
  assign _13007_ = \bapg_rd.w_ptr_r [3] ? _13006_ : _12999_;
  assign _13008_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [11] : \MSYNC_1r1w.synth.nz.mem[688] [11];
  assign _13009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [11] : \MSYNC_1r1w.synth.nz.mem[690] [11];
  assign _13010_ = \bapg_rd.w_ptr_r [1] ? _13009_ : _13008_;
  assign _13011_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [11] : \MSYNC_1r1w.synth.nz.mem[692] [11];
  assign _13012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [11] : \MSYNC_1r1w.synth.nz.mem[694] [11];
  assign _13013_ = \bapg_rd.w_ptr_r [1] ? _13012_ : _13011_;
  assign _13014_ = \bapg_rd.w_ptr_r [2] ? _13013_ : _13010_;
  assign _13015_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [11] : \MSYNC_1r1w.synth.nz.mem[696] [11];
  assign _13016_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [11] : \MSYNC_1r1w.synth.nz.mem[698] [11];
  assign _13017_ = \bapg_rd.w_ptr_r [1] ? _13016_ : _13015_;
  assign _13018_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [11] : \MSYNC_1r1w.synth.nz.mem[700] [11];
  assign _13019_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [11] : \MSYNC_1r1w.synth.nz.mem[702] [11];
  assign _13020_ = \bapg_rd.w_ptr_r [1] ? _13019_ : _13018_;
  assign _13021_ = \bapg_rd.w_ptr_r [2] ? _13020_ : _13017_;
  assign _13022_ = \bapg_rd.w_ptr_r [3] ? _13021_ : _13014_;
  assign _13023_ = \bapg_rd.w_ptr_r [4] ? _13022_ : _13007_;
  assign _13024_ = \bapg_rd.w_ptr_r [5] ? _13023_ : _12992_;
  assign _13025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [11] : \MSYNC_1r1w.synth.nz.mem[704] [11];
  assign _13026_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [11] : \MSYNC_1r1w.synth.nz.mem[706] [11];
  assign _13027_ = \bapg_rd.w_ptr_r [1] ? _13026_ : _13025_;
  assign _13028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [11] : \MSYNC_1r1w.synth.nz.mem[708] [11];
  assign _13029_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [11] : \MSYNC_1r1w.synth.nz.mem[710] [11];
  assign _13030_ = \bapg_rd.w_ptr_r [1] ? _13029_ : _13028_;
  assign _13031_ = \bapg_rd.w_ptr_r [2] ? _13030_ : _13027_;
  assign _13032_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [11] : \MSYNC_1r1w.synth.nz.mem[712] [11];
  assign _13033_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [11] : \MSYNC_1r1w.synth.nz.mem[714] [11];
  assign _13034_ = \bapg_rd.w_ptr_r [1] ? _13033_ : _13032_;
  assign _13035_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [11] : \MSYNC_1r1w.synth.nz.mem[716] [11];
  assign _13036_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [11] : \MSYNC_1r1w.synth.nz.mem[718] [11];
  assign _13037_ = \bapg_rd.w_ptr_r [1] ? _13036_ : _13035_;
  assign _13038_ = \bapg_rd.w_ptr_r [2] ? _13037_ : _13034_;
  assign _13039_ = \bapg_rd.w_ptr_r [3] ? _13038_ : _13031_;
  assign _13040_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [11] : \MSYNC_1r1w.synth.nz.mem[720] [11];
  assign _13041_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [11] : \MSYNC_1r1w.synth.nz.mem[722] [11];
  assign _13042_ = \bapg_rd.w_ptr_r [1] ? _13041_ : _13040_;
  assign _13043_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [11] : \MSYNC_1r1w.synth.nz.mem[724] [11];
  assign _13044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [11] : \MSYNC_1r1w.synth.nz.mem[726] [11];
  assign _13045_ = \bapg_rd.w_ptr_r [1] ? _13044_ : _13043_;
  assign _13046_ = \bapg_rd.w_ptr_r [2] ? _13045_ : _13042_;
  assign _13047_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [11] : \MSYNC_1r1w.synth.nz.mem[728] [11];
  assign _13048_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [11] : \MSYNC_1r1w.synth.nz.mem[730] [11];
  assign _13049_ = \bapg_rd.w_ptr_r [1] ? _13048_ : _13047_;
  assign _13050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [11] : \MSYNC_1r1w.synth.nz.mem[732] [11];
  assign _13051_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [11] : \MSYNC_1r1w.synth.nz.mem[734] [11];
  assign _13052_ = \bapg_rd.w_ptr_r [1] ? _13051_ : _13050_;
  assign _13053_ = \bapg_rd.w_ptr_r [2] ? _13052_ : _13049_;
  assign _13054_ = \bapg_rd.w_ptr_r [3] ? _13053_ : _13046_;
  assign _13055_ = \bapg_rd.w_ptr_r [4] ? _13054_ : _13039_;
  assign _13056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [11] : \MSYNC_1r1w.synth.nz.mem[736] [11];
  assign _13057_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [11] : \MSYNC_1r1w.synth.nz.mem[738] [11];
  assign _13058_ = \bapg_rd.w_ptr_r [1] ? _13057_ : _13056_;
  assign _13059_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [11] : \MSYNC_1r1w.synth.nz.mem[740] [11];
  assign _13060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [11] : \MSYNC_1r1w.synth.nz.mem[742] [11];
  assign _13061_ = \bapg_rd.w_ptr_r [1] ? _13060_ : _13059_;
  assign _13062_ = \bapg_rd.w_ptr_r [2] ? _13061_ : _13058_;
  assign _13063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [11] : \MSYNC_1r1w.synth.nz.mem[744] [11];
  assign _13064_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [11] : \MSYNC_1r1w.synth.nz.mem[746] [11];
  assign _13065_ = \bapg_rd.w_ptr_r [1] ? _13064_ : _13063_;
  assign _13066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [11] : \MSYNC_1r1w.synth.nz.mem[748] [11];
  assign _13067_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [11] : \MSYNC_1r1w.synth.nz.mem[750] [11];
  assign _13068_ = \bapg_rd.w_ptr_r [1] ? _13067_ : _13066_;
  assign _13069_ = \bapg_rd.w_ptr_r [2] ? _13068_ : _13065_;
  assign _13070_ = \bapg_rd.w_ptr_r [3] ? _13069_ : _13062_;
  assign _13071_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [11] : \MSYNC_1r1w.synth.nz.mem[752] [11];
  assign _13072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [11] : \MSYNC_1r1w.synth.nz.mem[754] [11];
  assign _13073_ = \bapg_rd.w_ptr_r [1] ? _13072_ : _13071_;
  assign _13074_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [11] : \MSYNC_1r1w.synth.nz.mem[756] [11];
  assign _13075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [11] : \MSYNC_1r1w.synth.nz.mem[758] [11];
  assign _13076_ = \bapg_rd.w_ptr_r [1] ? _13075_ : _13074_;
  assign _13077_ = \bapg_rd.w_ptr_r [2] ? _13076_ : _13073_;
  assign _13078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [11] : \MSYNC_1r1w.synth.nz.mem[760] [11];
  assign _13079_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [11] : \MSYNC_1r1w.synth.nz.mem[762] [11];
  assign _13080_ = \bapg_rd.w_ptr_r [1] ? _13079_ : _13078_;
  assign _13081_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [11] : \MSYNC_1r1w.synth.nz.mem[764] [11];
  assign _13082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [11] : \MSYNC_1r1w.synth.nz.mem[766] [11];
  assign _13083_ = \bapg_rd.w_ptr_r [1] ? _13082_ : _13081_;
  assign _13084_ = \bapg_rd.w_ptr_r [2] ? _13083_ : _13080_;
  assign _13085_ = \bapg_rd.w_ptr_r [3] ? _13084_ : _13077_;
  assign _13086_ = \bapg_rd.w_ptr_r [4] ? _13085_ : _13070_;
  assign _13087_ = \bapg_rd.w_ptr_r [5] ? _13086_ : _13055_;
  assign _13088_ = \bapg_rd.w_ptr_r [6] ? _13087_ : _13024_;
  assign _13089_ = \bapg_rd.w_ptr_r [7] ? _13088_ : _12961_;
  assign _13090_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [11] : \MSYNC_1r1w.synth.nz.mem[768] [11];
  assign _13091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [11] : \MSYNC_1r1w.synth.nz.mem[770] [11];
  assign _13092_ = \bapg_rd.w_ptr_r [1] ? _13091_ : _13090_;
  assign _13093_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [11] : \MSYNC_1r1w.synth.nz.mem[772] [11];
  assign _13094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [11] : \MSYNC_1r1w.synth.nz.mem[774] [11];
  assign _13095_ = \bapg_rd.w_ptr_r [1] ? _13094_ : _13093_;
  assign _13096_ = \bapg_rd.w_ptr_r [2] ? _13095_ : _13092_;
  assign _13097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [11] : \MSYNC_1r1w.synth.nz.mem[776] [11];
  assign _13098_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [11] : \MSYNC_1r1w.synth.nz.mem[778] [11];
  assign _13099_ = \bapg_rd.w_ptr_r [1] ? _13098_ : _13097_;
  assign _13100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [11] : \MSYNC_1r1w.synth.nz.mem[780] [11];
  assign _13101_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [11] : \MSYNC_1r1w.synth.nz.mem[782] [11];
  assign _13102_ = \bapg_rd.w_ptr_r [1] ? _13101_ : _13100_;
  assign _13103_ = \bapg_rd.w_ptr_r [2] ? _13102_ : _13099_;
  assign _13104_ = \bapg_rd.w_ptr_r [3] ? _13103_ : _13096_;
  assign _13105_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [11] : \MSYNC_1r1w.synth.nz.mem[784] [11];
  assign _13106_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [11] : \MSYNC_1r1w.synth.nz.mem[786] [11];
  assign _13107_ = \bapg_rd.w_ptr_r [1] ? _13106_ : _13105_;
  assign _13108_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [11] : \MSYNC_1r1w.synth.nz.mem[788] [11];
  assign _13109_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [11] : \MSYNC_1r1w.synth.nz.mem[790] [11];
  assign _13110_ = \bapg_rd.w_ptr_r [1] ? _13109_ : _13108_;
  assign _13111_ = \bapg_rd.w_ptr_r [2] ? _13110_ : _13107_;
  assign _13112_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [11] : \MSYNC_1r1w.synth.nz.mem[792] [11];
  assign _13113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [11] : \MSYNC_1r1w.synth.nz.mem[794] [11];
  assign _13114_ = \bapg_rd.w_ptr_r [1] ? _13113_ : _13112_;
  assign _13115_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [11] : \MSYNC_1r1w.synth.nz.mem[796] [11];
  assign _13116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [11] : \MSYNC_1r1w.synth.nz.mem[798] [11];
  assign _13117_ = \bapg_rd.w_ptr_r [1] ? _13116_ : _13115_;
  assign _13118_ = \bapg_rd.w_ptr_r [2] ? _13117_ : _13114_;
  assign _13119_ = \bapg_rd.w_ptr_r [3] ? _13118_ : _13111_;
  assign _13120_ = \bapg_rd.w_ptr_r [4] ? _13119_ : _13104_;
  assign _13121_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [11] : \MSYNC_1r1w.synth.nz.mem[800] [11];
  assign _13122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [11] : \MSYNC_1r1w.synth.nz.mem[802] [11];
  assign _13123_ = \bapg_rd.w_ptr_r [1] ? _13122_ : _13121_;
  assign _13124_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [11] : \MSYNC_1r1w.synth.nz.mem[804] [11];
  assign _13125_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [11] : \MSYNC_1r1w.synth.nz.mem[806] [11];
  assign _13126_ = \bapg_rd.w_ptr_r [1] ? _13125_ : _13124_;
  assign _13127_ = \bapg_rd.w_ptr_r [2] ? _13126_ : _13123_;
  assign _13128_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [11] : \MSYNC_1r1w.synth.nz.mem[808] [11];
  assign _13129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [11] : \MSYNC_1r1w.synth.nz.mem[810] [11];
  assign _13130_ = \bapg_rd.w_ptr_r [1] ? _13129_ : _13128_;
  assign _13131_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [11] : \MSYNC_1r1w.synth.nz.mem[812] [11];
  assign _13132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [11] : \MSYNC_1r1w.synth.nz.mem[814] [11];
  assign _13133_ = \bapg_rd.w_ptr_r [1] ? _13132_ : _13131_;
  assign _13134_ = \bapg_rd.w_ptr_r [2] ? _13133_ : _13130_;
  assign _13135_ = \bapg_rd.w_ptr_r [3] ? _13134_ : _13127_;
  assign _13136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [11] : \MSYNC_1r1w.synth.nz.mem[816] [11];
  assign _13137_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [11] : \MSYNC_1r1w.synth.nz.mem[818] [11];
  assign _13138_ = \bapg_rd.w_ptr_r [1] ? _13137_ : _13136_;
  assign _13139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [11] : \MSYNC_1r1w.synth.nz.mem[820] [11];
  assign _13140_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [11] : \MSYNC_1r1w.synth.nz.mem[822] [11];
  assign _13141_ = \bapg_rd.w_ptr_r [1] ? _13140_ : _13139_;
  assign _13142_ = \bapg_rd.w_ptr_r [2] ? _13141_ : _13138_;
  assign _13143_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [11] : \MSYNC_1r1w.synth.nz.mem[824] [11];
  assign _13144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [11] : \MSYNC_1r1w.synth.nz.mem[826] [11];
  assign _13145_ = \bapg_rd.w_ptr_r [1] ? _13144_ : _13143_;
  assign _13146_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [11] : \MSYNC_1r1w.synth.nz.mem[828] [11];
  assign _13147_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [11] : \MSYNC_1r1w.synth.nz.mem[830] [11];
  assign _13148_ = \bapg_rd.w_ptr_r [1] ? _13147_ : _13146_;
  assign _13149_ = \bapg_rd.w_ptr_r [2] ? _13148_ : _13145_;
  assign _13150_ = \bapg_rd.w_ptr_r [3] ? _13149_ : _13142_;
  assign _13151_ = \bapg_rd.w_ptr_r [4] ? _13150_ : _13135_;
  assign _13152_ = \bapg_rd.w_ptr_r [5] ? _13151_ : _13120_;
  assign _13153_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [11] : \MSYNC_1r1w.synth.nz.mem[832] [11];
  assign _13154_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [11] : \MSYNC_1r1w.synth.nz.mem[834] [11];
  assign _13155_ = \bapg_rd.w_ptr_r [1] ? _13154_ : _13153_;
  assign _13156_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [11] : \MSYNC_1r1w.synth.nz.mem[836] [11];
  assign _13157_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [11] : \MSYNC_1r1w.synth.nz.mem[838] [11];
  assign _13158_ = \bapg_rd.w_ptr_r [1] ? _13157_ : _13156_;
  assign _13159_ = \bapg_rd.w_ptr_r [2] ? _13158_ : _13155_;
  assign _13160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [11] : \MSYNC_1r1w.synth.nz.mem[840] [11];
  assign _13161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [11] : \MSYNC_1r1w.synth.nz.mem[842] [11];
  assign _13162_ = \bapg_rd.w_ptr_r [1] ? _13161_ : _13160_;
  assign _13163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [11] : \MSYNC_1r1w.synth.nz.mem[844] [11];
  assign _13164_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [11] : \MSYNC_1r1w.synth.nz.mem[846] [11];
  assign _13165_ = \bapg_rd.w_ptr_r [1] ? _13164_ : _13163_;
  assign _13166_ = \bapg_rd.w_ptr_r [2] ? _13165_ : _13162_;
  assign _13167_ = \bapg_rd.w_ptr_r [3] ? _13166_ : _13159_;
  assign _13168_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [11] : \MSYNC_1r1w.synth.nz.mem[848] [11];
  assign _13169_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [11] : \MSYNC_1r1w.synth.nz.mem[850] [11];
  assign _13170_ = \bapg_rd.w_ptr_r [1] ? _13169_ : _13168_;
  assign _13171_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [11] : \MSYNC_1r1w.synth.nz.mem[852] [11];
  assign _13172_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [11] : \MSYNC_1r1w.synth.nz.mem[854] [11];
  assign _13173_ = \bapg_rd.w_ptr_r [1] ? _13172_ : _13171_;
  assign _13174_ = \bapg_rd.w_ptr_r [2] ? _13173_ : _13170_;
  assign _13175_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [11] : \MSYNC_1r1w.synth.nz.mem[856] [11];
  assign _13176_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [11] : \MSYNC_1r1w.synth.nz.mem[858] [11];
  assign _13177_ = \bapg_rd.w_ptr_r [1] ? _13176_ : _13175_;
  assign _13178_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [11] : \MSYNC_1r1w.synth.nz.mem[860] [11];
  assign _13179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [11] : \MSYNC_1r1w.synth.nz.mem[862] [11];
  assign _13180_ = \bapg_rd.w_ptr_r [1] ? _13179_ : _13178_;
  assign _13181_ = \bapg_rd.w_ptr_r [2] ? _13180_ : _13177_;
  assign _13182_ = \bapg_rd.w_ptr_r [3] ? _13181_ : _13174_;
  assign _13183_ = \bapg_rd.w_ptr_r [4] ? _13182_ : _13167_;
  assign _13184_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [11] : \MSYNC_1r1w.synth.nz.mem[864] [11];
  assign _13185_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [11] : \MSYNC_1r1w.synth.nz.mem[866] [11];
  assign _13186_ = \bapg_rd.w_ptr_r [1] ? _13185_ : _13184_;
  assign _13187_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [11] : \MSYNC_1r1w.synth.nz.mem[868] [11];
  assign _13188_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [11] : \MSYNC_1r1w.synth.nz.mem[870] [11];
  assign _13189_ = \bapg_rd.w_ptr_r [1] ? _13188_ : _13187_;
  assign _13190_ = \bapg_rd.w_ptr_r [2] ? _13189_ : _13186_;
  assign _13191_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [11] : \MSYNC_1r1w.synth.nz.mem[872] [11];
  assign _13192_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [11] : \MSYNC_1r1w.synth.nz.mem[874] [11];
  assign _13193_ = \bapg_rd.w_ptr_r [1] ? _13192_ : _13191_;
  assign _13194_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [11] : \MSYNC_1r1w.synth.nz.mem[876] [11];
  assign _13195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [11] : \MSYNC_1r1w.synth.nz.mem[878] [11];
  assign _13196_ = \bapg_rd.w_ptr_r [1] ? _13195_ : _13194_;
  assign _13197_ = \bapg_rd.w_ptr_r [2] ? _13196_ : _13193_;
  assign _13198_ = \bapg_rd.w_ptr_r [3] ? _13197_ : _13190_;
  assign _13199_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [11] : \MSYNC_1r1w.synth.nz.mem[880] [11];
  assign _13200_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [11] : \MSYNC_1r1w.synth.nz.mem[882] [11];
  assign _13201_ = \bapg_rd.w_ptr_r [1] ? _13200_ : _13199_;
  assign _13202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [11] : \MSYNC_1r1w.synth.nz.mem[884] [11];
  assign _13203_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [11] : \MSYNC_1r1w.synth.nz.mem[886] [11];
  assign _13204_ = \bapg_rd.w_ptr_r [1] ? _13203_ : _13202_;
  assign _13205_ = \bapg_rd.w_ptr_r [2] ? _13204_ : _13201_;
  assign _13206_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [11] : \MSYNC_1r1w.synth.nz.mem[888] [11];
  assign _13207_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [11] : \MSYNC_1r1w.synth.nz.mem[890] [11];
  assign _13208_ = \bapg_rd.w_ptr_r [1] ? _13207_ : _13206_;
  assign _13209_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [11] : \MSYNC_1r1w.synth.nz.mem[892] [11];
  assign _13210_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [11] : \MSYNC_1r1w.synth.nz.mem[894] [11];
  assign _13211_ = \bapg_rd.w_ptr_r [1] ? _13210_ : _13209_;
  assign _13212_ = \bapg_rd.w_ptr_r [2] ? _13211_ : _13208_;
  assign _13213_ = \bapg_rd.w_ptr_r [3] ? _13212_ : _13205_;
  assign _13214_ = \bapg_rd.w_ptr_r [4] ? _13213_ : _13198_;
  assign _13215_ = \bapg_rd.w_ptr_r [5] ? _13214_ : _13183_;
  assign _13216_ = \bapg_rd.w_ptr_r [6] ? _13215_ : _13152_;
  assign _13217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [11] : \MSYNC_1r1w.synth.nz.mem[896] [11];
  assign _13218_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [11] : \MSYNC_1r1w.synth.nz.mem[898] [11];
  assign _13219_ = \bapg_rd.w_ptr_r [1] ? _13218_ : _13217_;
  assign _13220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [11] : \MSYNC_1r1w.synth.nz.mem[900] [11];
  assign _13221_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [11] : \MSYNC_1r1w.synth.nz.mem[902] [11];
  assign _13222_ = \bapg_rd.w_ptr_r [1] ? _13221_ : _13220_;
  assign _13223_ = \bapg_rd.w_ptr_r [2] ? _13222_ : _13219_;
  assign _13224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [11] : \MSYNC_1r1w.synth.nz.mem[904] [11];
  assign _13225_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [11] : \MSYNC_1r1w.synth.nz.mem[906] [11];
  assign _13226_ = \bapg_rd.w_ptr_r [1] ? _13225_ : _13224_;
  assign _13227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [11] : \MSYNC_1r1w.synth.nz.mem[908] [11];
  assign _13228_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [11] : \MSYNC_1r1w.synth.nz.mem[910] [11];
  assign _13229_ = \bapg_rd.w_ptr_r [1] ? _13228_ : _13227_;
  assign _13230_ = \bapg_rd.w_ptr_r [2] ? _13229_ : _13226_;
  assign _13231_ = \bapg_rd.w_ptr_r [3] ? _13230_ : _13223_;
  assign _13232_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [11] : \MSYNC_1r1w.synth.nz.mem[912] [11];
  assign _13233_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [11] : \MSYNC_1r1w.synth.nz.mem[914] [11];
  assign _13234_ = \bapg_rd.w_ptr_r [1] ? _13233_ : _13232_;
  assign _13235_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [11] : \MSYNC_1r1w.synth.nz.mem[916] [11];
  assign _13236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [11] : \MSYNC_1r1w.synth.nz.mem[918] [11];
  assign _13237_ = \bapg_rd.w_ptr_r [1] ? _13236_ : _13235_;
  assign _13238_ = \bapg_rd.w_ptr_r [2] ? _13237_ : _13234_;
  assign _13239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [11] : \MSYNC_1r1w.synth.nz.mem[920] [11];
  assign _13240_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [11] : \MSYNC_1r1w.synth.nz.mem[922] [11];
  assign _13241_ = \bapg_rd.w_ptr_r [1] ? _13240_ : _13239_;
  assign _13242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [11] : \MSYNC_1r1w.synth.nz.mem[924] [11];
  assign _13243_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [11] : \MSYNC_1r1w.synth.nz.mem[926] [11];
  assign _13244_ = \bapg_rd.w_ptr_r [1] ? _13243_ : _13242_;
  assign _13245_ = \bapg_rd.w_ptr_r [2] ? _13244_ : _13241_;
  assign _13246_ = \bapg_rd.w_ptr_r [3] ? _13245_ : _13238_;
  assign _13247_ = \bapg_rd.w_ptr_r [4] ? _13246_ : _13231_;
  assign _13248_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [11] : \MSYNC_1r1w.synth.nz.mem[928] [11];
  assign _13249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [11] : \MSYNC_1r1w.synth.nz.mem[930] [11];
  assign _13250_ = \bapg_rd.w_ptr_r [1] ? _13249_ : _13248_;
  assign _13251_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [11] : \MSYNC_1r1w.synth.nz.mem[932] [11];
  assign _13252_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [11] : \MSYNC_1r1w.synth.nz.mem[934] [11];
  assign _13253_ = \bapg_rd.w_ptr_r [1] ? _13252_ : _13251_;
  assign _13254_ = \bapg_rd.w_ptr_r [2] ? _13253_ : _13250_;
  assign _13255_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [11] : \MSYNC_1r1w.synth.nz.mem[936] [11];
  assign _13256_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [11] : \MSYNC_1r1w.synth.nz.mem[938] [11];
  assign _13257_ = \bapg_rd.w_ptr_r [1] ? _13256_ : _13255_;
  assign _13258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [11] : \MSYNC_1r1w.synth.nz.mem[940] [11];
  assign _13259_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [11] : \MSYNC_1r1w.synth.nz.mem[942] [11];
  assign _13260_ = \bapg_rd.w_ptr_r [1] ? _13259_ : _13258_;
  assign _13261_ = \bapg_rd.w_ptr_r [2] ? _13260_ : _13257_;
  assign _13262_ = \bapg_rd.w_ptr_r [3] ? _13261_ : _13254_;
  assign _13263_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [11] : \MSYNC_1r1w.synth.nz.mem[944] [11];
  assign _13264_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [11] : \MSYNC_1r1w.synth.nz.mem[946] [11];
  assign _13265_ = \bapg_rd.w_ptr_r [1] ? _13264_ : _13263_;
  assign _13266_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [11] : \MSYNC_1r1w.synth.nz.mem[948] [11];
  assign _13267_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [11] : \MSYNC_1r1w.synth.nz.mem[950] [11];
  assign _13268_ = \bapg_rd.w_ptr_r [1] ? _13267_ : _13266_;
  assign _13269_ = \bapg_rd.w_ptr_r [2] ? _13268_ : _13265_;
  assign _13270_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [11] : \MSYNC_1r1w.synth.nz.mem[952] [11];
  assign _13271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [11] : \MSYNC_1r1w.synth.nz.mem[954] [11];
  assign _13272_ = \bapg_rd.w_ptr_r [1] ? _13271_ : _13270_;
  assign _13273_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [11] : \MSYNC_1r1w.synth.nz.mem[956] [11];
  assign _13274_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [11] : \MSYNC_1r1w.synth.nz.mem[958] [11];
  assign _13275_ = \bapg_rd.w_ptr_r [1] ? _13274_ : _13273_;
  assign _13276_ = \bapg_rd.w_ptr_r [2] ? _13275_ : _13272_;
  assign _13277_ = \bapg_rd.w_ptr_r [3] ? _13276_ : _13269_;
  assign _13278_ = \bapg_rd.w_ptr_r [4] ? _13277_ : _13262_;
  assign _13279_ = \bapg_rd.w_ptr_r [5] ? _13278_ : _13247_;
  assign _13280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [11] : \MSYNC_1r1w.synth.nz.mem[960] [11];
  assign _13281_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [11] : \MSYNC_1r1w.synth.nz.mem[962] [11];
  assign _13282_ = \bapg_rd.w_ptr_r [1] ? _13281_ : _13280_;
  assign _13283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [11] : \MSYNC_1r1w.synth.nz.mem[964] [11];
  assign _13284_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [11] : \MSYNC_1r1w.synth.nz.mem[966] [11];
  assign _13285_ = \bapg_rd.w_ptr_r [1] ? _13284_ : _13283_;
  assign _13286_ = \bapg_rd.w_ptr_r [2] ? _13285_ : _13282_;
  assign _13287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [11] : \MSYNC_1r1w.synth.nz.mem[968] [11];
  assign _13288_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [11] : \MSYNC_1r1w.synth.nz.mem[970] [11];
  assign _13289_ = \bapg_rd.w_ptr_r [1] ? _13288_ : _13287_;
  assign _13290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [11] : \MSYNC_1r1w.synth.nz.mem[972] [11];
  assign _13291_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [11] : \MSYNC_1r1w.synth.nz.mem[974] [11];
  assign _13292_ = \bapg_rd.w_ptr_r [1] ? _13291_ : _13290_;
  assign _13293_ = \bapg_rd.w_ptr_r [2] ? _13292_ : _13289_;
  assign _13294_ = \bapg_rd.w_ptr_r [3] ? _13293_ : _13286_;
  assign _13295_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [11] : \MSYNC_1r1w.synth.nz.mem[976] [11];
  assign _13296_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [11] : \MSYNC_1r1w.synth.nz.mem[978] [11];
  assign _13297_ = \bapg_rd.w_ptr_r [1] ? _13296_ : _13295_;
  assign _13298_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [11] : \MSYNC_1r1w.synth.nz.mem[980] [11];
  assign _13299_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [11] : \MSYNC_1r1w.synth.nz.mem[982] [11];
  assign _13300_ = \bapg_rd.w_ptr_r [1] ? _13299_ : _13298_;
  assign _13301_ = \bapg_rd.w_ptr_r [2] ? _13300_ : _13297_;
  assign _13302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [11] : \MSYNC_1r1w.synth.nz.mem[984] [11];
  assign _13303_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [11] : \MSYNC_1r1w.synth.nz.mem[986] [11];
  assign _13304_ = \bapg_rd.w_ptr_r [1] ? _13303_ : _13302_;
  assign _13305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [11] : \MSYNC_1r1w.synth.nz.mem[988] [11];
  assign _13306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [11] : \MSYNC_1r1w.synth.nz.mem[990] [11];
  assign _13307_ = \bapg_rd.w_ptr_r [1] ? _13306_ : _13305_;
  assign _13308_ = \bapg_rd.w_ptr_r [2] ? _13307_ : _13304_;
  assign _13309_ = \bapg_rd.w_ptr_r [3] ? _13308_ : _13301_;
  assign _13310_ = \bapg_rd.w_ptr_r [4] ? _13309_ : _13294_;
  assign _13311_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [11] : \MSYNC_1r1w.synth.nz.mem[992] [11];
  assign _13312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [11] : \MSYNC_1r1w.synth.nz.mem[994] [11];
  assign _13313_ = \bapg_rd.w_ptr_r [1] ? _13312_ : _13311_;
  assign _13314_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [11] : \MSYNC_1r1w.synth.nz.mem[996] [11];
  assign _13315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [11] : \MSYNC_1r1w.synth.nz.mem[998] [11];
  assign _13316_ = \bapg_rd.w_ptr_r [1] ? _13315_ : _13314_;
  assign _13317_ = \bapg_rd.w_ptr_r [2] ? _13316_ : _13313_;
  assign _13318_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [11] : \MSYNC_1r1w.synth.nz.mem[1000] [11];
  assign _13319_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [11] : \MSYNC_1r1w.synth.nz.mem[1002] [11];
  assign _13320_ = \bapg_rd.w_ptr_r [1] ? _13319_ : _13318_;
  assign _13321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [11] : \MSYNC_1r1w.synth.nz.mem[1004] [11];
  assign _13322_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [11] : \MSYNC_1r1w.synth.nz.mem[1006] [11];
  assign _13323_ = \bapg_rd.w_ptr_r [1] ? _13322_ : _13321_;
  assign _13324_ = \bapg_rd.w_ptr_r [2] ? _13323_ : _13320_;
  assign _13325_ = \bapg_rd.w_ptr_r [3] ? _13324_ : _13317_;
  assign _13326_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [11] : \MSYNC_1r1w.synth.nz.mem[1008] [11];
  assign _13327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [11] : \MSYNC_1r1w.synth.nz.mem[1010] [11];
  assign _13328_ = \bapg_rd.w_ptr_r [1] ? _13327_ : _13326_;
  assign _13329_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [11] : \MSYNC_1r1w.synth.nz.mem[1012] [11];
  assign _13330_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [11] : \MSYNC_1r1w.synth.nz.mem[1014] [11];
  assign _13331_ = \bapg_rd.w_ptr_r [1] ? _13330_ : _13329_;
  assign _13332_ = \bapg_rd.w_ptr_r [2] ? _13331_ : _13328_;
  assign _13333_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [11] : \MSYNC_1r1w.synth.nz.mem[1016] [11];
  assign _13334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [11] : \MSYNC_1r1w.synth.nz.mem[1018] [11];
  assign _13335_ = \bapg_rd.w_ptr_r [1] ? _13334_ : _13333_;
  assign _13336_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [11] : \MSYNC_1r1w.synth.nz.mem[1020] [11];
  assign _13337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [11] : \MSYNC_1r1w.synth.nz.mem[1022] [11];
  assign _13338_ = \bapg_rd.w_ptr_r [1] ? _13337_ : _13336_;
  assign _13339_ = \bapg_rd.w_ptr_r [2] ? _13338_ : _13335_;
  assign _13340_ = \bapg_rd.w_ptr_r [3] ? _13339_ : _13332_;
  assign _13341_ = \bapg_rd.w_ptr_r [4] ? _13340_ : _13325_;
  assign _13342_ = \bapg_rd.w_ptr_r [5] ? _13341_ : _13310_;
  assign _13343_ = \bapg_rd.w_ptr_r [6] ? _13342_ : _13279_;
  assign _13344_ = \bapg_rd.w_ptr_r [7] ? _13343_ : _13216_;
  assign _13345_ = \bapg_rd.w_ptr_r [8] ? _13344_ : _13089_;
  assign r_data_o[11] = \bapg_rd.w_ptr_r [9] ? _13345_ : _12834_;
  assign _13346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [12] : \MSYNC_1r1w.synth.nz.mem[0] [12];
  assign _13347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [12] : \MSYNC_1r1w.synth.nz.mem[2] [12];
  assign _13348_ = \bapg_rd.w_ptr_r [1] ? _13347_ : _13346_;
  assign _13349_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [12] : \MSYNC_1r1w.synth.nz.mem[4] [12];
  assign _13350_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [12] : \MSYNC_1r1w.synth.nz.mem[6] [12];
  assign _13351_ = \bapg_rd.w_ptr_r [1] ? _13350_ : _13349_;
  assign _13352_ = \bapg_rd.w_ptr_r [2] ? _13351_ : _13348_;
  assign _13353_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [12] : \MSYNC_1r1w.synth.nz.mem[8] [12];
  assign _13354_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [12] : \MSYNC_1r1w.synth.nz.mem[10] [12];
  assign _13355_ = \bapg_rd.w_ptr_r [1] ? _13354_ : _13353_;
  assign _13356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [12] : \MSYNC_1r1w.synth.nz.mem[12] [12];
  assign _13357_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [12] : \MSYNC_1r1w.synth.nz.mem[14] [12];
  assign _13358_ = \bapg_rd.w_ptr_r [1] ? _13357_ : _13356_;
  assign _13359_ = \bapg_rd.w_ptr_r [2] ? _13358_ : _13355_;
  assign _13360_ = \bapg_rd.w_ptr_r [3] ? _13359_ : _13352_;
  assign _13361_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [12] : \MSYNC_1r1w.synth.nz.mem[16] [12];
  assign _13362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [12] : \MSYNC_1r1w.synth.nz.mem[18] [12];
  assign _13363_ = \bapg_rd.w_ptr_r [1] ? _13362_ : _13361_;
  assign _13364_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [12] : \MSYNC_1r1w.synth.nz.mem[20] [12];
  assign _13365_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [12] : \MSYNC_1r1w.synth.nz.mem[22] [12];
  assign _13366_ = \bapg_rd.w_ptr_r [1] ? _13365_ : _13364_;
  assign _13367_ = \bapg_rd.w_ptr_r [2] ? _13366_ : _13363_;
  assign _13368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [12] : \MSYNC_1r1w.synth.nz.mem[24] [12];
  assign _13369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [12] : \MSYNC_1r1w.synth.nz.mem[26] [12];
  assign _13370_ = \bapg_rd.w_ptr_r [1] ? _13369_ : _13368_;
  assign _13371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [12] : \MSYNC_1r1w.synth.nz.mem[28] [12];
  assign _13372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [12] : \MSYNC_1r1w.synth.nz.mem[30] [12];
  assign _13373_ = \bapg_rd.w_ptr_r [1] ? _13372_ : _13371_;
  assign _13374_ = \bapg_rd.w_ptr_r [2] ? _13373_ : _13370_;
  assign _13375_ = \bapg_rd.w_ptr_r [3] ? _13374_ : _13367_;
  assign _13376_ = \bapg_rd.w_ptr_r [4] ? _13375_ : _13360_;
  assign _13377_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [12] : \MSYNC_1r1w.synth.nz.mem[32] [12];
  assign _13378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [12] : \MSYNC_1r1w.synth.nz.mem[34] [12];
  assign _13379_ = \bapg_rd.w_ptr_r [1] ? _13378_ : _13377_;
  assign _13380_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [12] : \MSYNC_1r1w.synth.nz.mem[36] [12];
  assign _13381_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [12] : \MSYNC_1r1w.synth.nz.mem[38] [12];
  assign _13382_ = \bapg_rd.w_ptr_r [1] ? _13381_ : _13380_;
  assign _13383_ = \bapg_rd.w_ptr_r [2] ? _13382_ : _13379_;
  assign _13384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [12] : \MSYNC_1r1w.synth.nz.mem[40] [12];
  assign _13385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [12] : \MSYNC_1r1w.synth.nz.mem[42] [12];
  assign _13386_ = \bapg_rd.w_ptr_r [1] ? _13385_ : _13384_;
  assign _13387_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [12] : \MSYNC_1r1w.synth.nz.mem[44] [12];
  assign _13388_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [12] : \MSYNC_1r1w.synth.nz.mem[46] [12];
  assign _13389_ = \bapg_rd.w_ptr_r [1] ? _13388_ : _13387_;
  assign _13390_ = \bapg_rd.w_ptr_r [2] ? _13389_ : _13386_;
  assign _13391_ = \bapg_rd.w_ptr_r [3] ? _13390_ : _13383_;
  assign _13392_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [12] : \MSYNC_1r1w.synth.nz.mem[48] [12];
  assign _13393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [12] : \MSYNC_1r1w.synth.nz.mem[50] [12];
  assign _13394_ = \bapg_rd.w_ptr_r [1] ? _13393_ : _13392_;
  assign _13395_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [12] : \MSYNC_1r1w.synth.nz.mem[52] [12];
  assign _13396_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [12] : \MSYNC_1r1w.synth.nz.mem[54] [12];
  assign _13397_ = \bapg_rd.w_ptr_r [1] ? _13396_ : _13395_;
  assign _13398_ = \bapg_rd.w_ptr_r [2] ? _13397_ : _13394_;
  assign _13399_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [12] : \MSYNC_1r1w.synth.nz.mem[56] [12];
  assign _13400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [12] : \MSYNC_1r1w.synth.nz.mem[58] [12];
  assign _13401_ = \bapg_rd.w_ptr_r [1] ? _13400_ : _13399_;
  assign _13402_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [12] : \MSYNC_1r1w.synth.nz.mem[60] [12];
  assign _13403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [12] : \MSYNC_1r1w.synth.nz.mem[62] [12];
  assign _13404_ = \bapg_rd.w_ptr_r [1] ? _13403_ : _13402_;
  assign _13405_ = \bapg_rd.w_ptr_r [2] ? _13404_ : _13401_;
  assign _13406_ = \bapg_rd.w_ptr_r [3] ? _13405_ : _13398_;
  assign _13407_ = \bapg_rd.w_ptr_r [4] ? _13406_ : _13391_;
  assign _13408_ = \bapg_rd.w_ptr_r [5] ? _13407_ : _13376_;
  assign _13409_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [12] : \MSYNC_1r1w.synth.nz.mem[64] [12];
  assign _13410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [12] : \MSYNC_1r1w.synth.nz.mem[66] [12];
  assign _13411_ = \bapg_rd.w_ptr_r [1] ? _13410_ : _13409_;
  assign _13412_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [12] : \MSYNC_1r1w.synth.nz.mem[68] [12];
  assign _13413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [12] : \MSYNC_1r1w.synth.nz.mem[70] [12];
  assign _13414_ = \bapg_rd.w_ptr_r [1] ? _13413_ : _13412_;
  assign _13415_ = \bapg_rd.w_ptr_r [2] ? _13414_ : _13411_;
  assign _13416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [12] : \MSYNC_1r1w.synth.nz.mem[72] [12];
  assign _13417_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [12] : \MSYNC_1r1w.synth.nz.mem[74] [12];
  assign _13418_ = \bapg_rd.w_ptr_r [1] ? _13417_ : _13416_;
  assign _13419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [12] : \MSYNC_1r1w.synth.nz.mem[76] [12];
  assign _13420_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [12] : \MSYNC_1r1w.synth.nz.mem[78] [12];
  assign _13421_ = \bapg_rd.w_ptr_r [1] ? _13420_ : _13419_;
  assign _13422_ = \bapg_rd.w_ptr_r [2] ? _13421_ : _13418_;
  assign _13423_ = \bapg_rd.w_ptr_r [3] ? _13422_ : _13415_;
  assign _13424_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [12] : \MSYNC_1r1w.synth.nz.mem[80] [12];
  assign _13425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [12] : \MSYNC_1r1w.synth.nz.mem[82] [12];
  assign _13426_ = \bapg_rd.w_ptr_r [1] ? _13425_ : _13424_;
  assign _13427_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [12] : \MSYNC_1r1w.synth.nz.mem[84] [12];
  assign _13428_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [12] : \MSYNC_1r1w.synth.nz.mem[86] [12];
  assign _13429_ = \bapg_rd.w_ptr_r [1] ? _13428_ : _13427_;
  assign _13430_ = \bapg_rd.w_ptr_r [2] ? _13429_ : _13426_;
  assign _13431_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [12] : \MSYNC_1r1w.synth.nz.mem[88] [12];
  assign _13432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [12] : \MSYNC_1r1w.synth.nz.mem[90] [12];
  assign _13433_ = \bapg_rd.w_ptr_r [1] ? _13432_ : _13431_;
  assign _13434_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [12] : \MSYNC_1r1w.synth.nz.mem[92] [12];
  assign _13435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [12] : \MSYNC_1r1w.synth.nz.mem[94] [12];
  assign _13436_ = \bapg_rd.w_ptr_r [1] ? _13435_ : _13434_;
  assign _13437_ = \bapg_rd.w_ptr_r [2] ? _13436_ : _13433_;
  assign _13438_ = \bapg_rd.w_ptr_r [3] ? _13437_ : _13430_;
  assign _13439_ = \bapg_rd.w_ptr_r [4] ? _13438_ : _13423_;
  assign _13440_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [12] : \MSYNC_1r1w.synth.nz.mem[96] [12];
  assign _13441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [12] : \MSYNC_1r1w.synth.nz.mem[98] [12];
  assign _13442_ = \bapg_rd.w_ptr_r [1] ? _13441_ : _13440_;
  assign _13443_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [12] : \MSYNC_1r1w.synth.nz.mem[100] [12];
  assign _13444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [12] : \MSYNC_1r1w.synth.nz.mem[102] [12];
  assign _13445_ = \bapg_rd.w_ptr_r [1] ? _13444_ : _13443_;
  assign _13446_ = \bapg_rd.w_ptr_r [2] ? _13445_ : _13442_;
  assign _13447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [12] : \MSYNC_1r1w.synth.nz.mem[104] [12];
  assign _13448_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [12] : \MSYNC_1r1w.synth.nz.mem[106] [12];
  assign _13449_ = \bapg_rd.w_ptr_r [1] ? _13448_ : _13447_;
  assign _13450_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [12] : \MSYNC_1r1w.synth.nz.mem[108] [12];
  assign _13451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [12] : \MSYNC_1r1w.synth.nz.mem[110] [12];
  assign _13452_ = \bapg_rd.w_ptr_r [1] ? _13451_ : _13450_;
  assign _13453_ = \bapg_rd.w_ptr_r [2] ? _13452_ : _13449_;
  assign _13454_ = \bapg_rd.w_ptr_r [3] ? _13453_ : _13446_;
  assign _13455_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [12] : \MSYNC_1r1w.synth.nz.mem[112] [12];
  assign _13456_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [12] : \MSYNC_1r1w.synth.nz.mem[114] [12];
  assign _13457_ = \bapg_rd.w_ptr_r [1] ? _13456_ : _13455_;
  assign _13458_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [12] : \MSYNC_1r1w.synth.nz.mem[116] [12];
  assign _13459_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [12] : \MSYNC_1r1w.synth.nz.mem[118] [12];
  assign _13460_ = \bapg_rd.w_ptr_r [1] ? _13459_ : _13458_;
  assign _13461_ = \bapg_rd.w_ptr_r [2] ? _13460_ : _13457_;
  assign _13462_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [12] : \MSYNC_1r1w.synth.nz.mem[120] [12];
  assign _13463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [12] : \MSYNC_1r1w.synth.nz.mem[122] [12];
  assign _13464_ = \bapg_rd.w_ptr_r [1] ? _13463_ : _13462_;
  assign _13465_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [12] : \MSYNC_1r1w.synth.nz.mem[124] [12];
  assign _13466_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [12] : \MSYNC_1r1w.synth.nz.mem[126] [12];
  assign _13467_ = \bapg_rd.w_ptr_r [1] ? _13466_ : _13465_;
  assign _13468_ = \bapg_rd.w_ptr_r [2] ? _13467_ : _13464_;
  assign _13469_ = \bapg_rd.w_ptr_r [3] ? _13468_ : _13461_;
  assign _13470_ = \bapg_rd.w_ptr_r [4] ? _13469_ : _13454_;
  assign _13471_ = \bapg_rd.w_ptr_r [5] ? _13470_ : _13439_;
  assign _13472_ = \bapg_rd.w_ptr_r [6] ? _13471_ : _13408_;
  assign _13473_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [12] : \MSYNC_1r1w.synth.nz.mem[128] [12];
  assign _13474_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [12] : \MSYNC_1r1w.synth.nz.mem[130] [12];
  assign _13475_ = \bapg_rd.w_ptr_r [1] ? _13474_ : _13473_;
  assign _13476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [12] : \MSYNC_1r1w.synth.nz.mem[132] [12];
  assign _13477_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [12] : \MSYNC_1r1w.synth.nz.mem[134] [12];
  assign _13478_ = \bapg_rd.w_ptr_r [1] ? _13477_ : _13476_;
  assign _13479_ = \bapg_rd.w_ptr_r [2] ? _13478_ : _13475_;
  assign _13480_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [12] : \MSYNC_1r1w.synth.nz.mem[136] [12];
  assign _13481_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [12] : \MSYNC_1r1w.synth.nz.mem[138] [12];
  assign _13482_ = \bapg_rd.w_ptr_r [1] ? _13481_ : _13480_;
  assign _13483_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [12] : \MSYNC_1r1w.synth.nz.mem[140] [12];
  assign _13484_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [12] : \MSYNC_1r1w.synth.nz.mem[142] [12];
  assign _13485_ = \bapg_rd.w_ptr_r [1] ? _13484_ : _13483_;
  assign _13486_ = \bapg_rd.w_ptr_r [2] ? _13485_ : _13482_;
  assign _13487_ = \bapg_rd.w_ptr_r [3] ? _13486_ : _13479_;
  assign _13488_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [12] : \MSYNC_1r1w.synth.nz.mem[144] [12];
  assign _13489_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [12] : \MSYNC_1r1w.synth.nz.mem[146] [12];
  assign _13490_ = \bapg_rd.w_ptr_r [1] ? _13489_ : _13488_;
  assign _13491_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [12] : \MSYNC_1r1w.synth.nz.mem[148] [12];
  assign _13492_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [12] : \MSYNC_1r1w.synth.nz.mem[150] [12];
  assign _13493_ = \bapg_rd.w_ptr_r [1] ? _13492_ : _13491_;
  assign _13494_ = \bapg_rd.w_ptr_r [2] ? _13493_ : _13490_;
  assign _13495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [12] : \MSYNC_1r1w.synth.nz.mem[152] [12];
  assign _13496_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [12] : \MSYNC_1r1w.synth.nz.mem[154] [12];
  assign _13497_ = \bapg_rd.w_ptr_r [1] ? _13496_ : _13495_;
  assign _13498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [12] : \MSYNC_1r1w.synth.nz.mem[156] [12];
  assign _13499_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [12] : \MSYNC_1r1w.synth.nz.mem[158] [12];
  assign _13500_ = \bapg_rd.w_ptr_r [1] ? _13499_ : _13498_;
  assign _13501_ = \bapg_rd.w_ptr_r [2] ? _13500_ : _13497_;
  assign _13502_ = \bapg_rd.w_ptr_r [3] ? _13501_ : _13494_;
  assign _13503_ = \bapg_rd.w_ptr_r [4] ? _13502_ : _13487_;
  assign _13504_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [12] : \MSYNC_1r1w.synth.nz.mem[160] [12];
  assign _13505_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [12] : \MSYNC_1r1w.synth.nz.mem[162] [12];
  assign _13506_ = \bapg_rd.w_ptr_r [1] ? _13505_ : _13504_;
  assign _13507_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [12] : \MSYNC_1r1w.synth.nz.mem[164] [12];
  assign _13508_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [12] : \MSYNC_1r1w.synth.nz.mem[166] [12];
  assign _13509_ = \bapg_rd.w_ptr_r [1] ? _13508_ : _13507_;
  assign _13510_ = \bapg_rd.w_ptr_r [2] ? _13509_ : _13506_;
  assign _13511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [12] : \MSYNC_1r1w.synth.nz.mem[168] [12];
  assign _13512_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [12] : \MSYNC_1r1w.synth.nz.mem[170] [12];
  assign _13513_ = \bapg_rd.w_ptr_r [1] ? _13512_ : _13511_;
  assign _13514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [12] : \MSYNC_1r1w.synth.nz.mem[172] [12];
  assign _13515_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [12] : \MSYNC_1r1w.synth.nz.mem[174] [12];
  assign _13516_ = \bapg_rd.w_ptr_r [1] ? _13515_ : _13514_;
  assign _13517_ = \bapg_rd.w_ptr_r [2] ? _13516_ : _13513_;
  assign _13518_ = \bapg_rd.w_ptr_r [3] ? _13517_ : _13510_;
  assign _13519_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [12] : \MSYNC_1r1w.synth.nz.mem[176] [12];
  assign _13520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [12] : \MSYNC_1r1w.synth.nz.mem[178] [12];
  assign _13521_ = \bapg_rd.w_ptr_r [1] ? _13520_ : _13519_;
  assign _13522_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [12] : \MSYNC_1r1w.synth.nz.mem[180] [12];
  assign _13523_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [12] : \MSYNC_1r1w.synth.nz.mem[182] [12];
  assign _13524_ = \bapg_rd.w_ptr_r [1] ? _13523_ : _13522_;
  assign _13525_ = \bapg_rd.w_ptr_r [2] ? _13524_ : _13521_;
  assign _13526_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [12] : \MSYNC_1r1w.synth.nz.mem[184] [12];
  assign _13527_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [12] : \MSYNC_1r1w.synth.nz.mem[186] [12];
  assign _13528_ = \bapg_rd.w_ptr_r [1] ? _13527_ : _13526_;
  assign _13529_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [12] : \MSYNC_1r1w.synth.nz.mem[188] [12];
  assign _13530_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [12] : \MSYNC_1r1w.synth.nz.mem[190] [12];
  assign _13531_ = \bapg_rd.w_ptr_r [1] ? _13530_ : _13529_;
  assign _13532_ = \bapg_rd.w_ptr_r [2] ? _13531_ : _13528_;
  assign _13533_ = \bapg_rd.w_ptr_r [3] ? _13532_ : _13525_;
  assign _13534_ = \bapg_rd.w_ptr_r [4] ? _13533_ : _13518_;
  assign _13535_ = \bapg_rd.w_ptr_r [5] ? _13534_ : _13503_;
  assign _13536_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [12] : \MSYNC_1r1w.synth.nz.mem[192] [12];
  assign _13537_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [12] : \MSYNC_1r1w.synth.nz.mem[194] [12];
  assign _13538_ = \bapg_rd.w_ptr_r [1] ? _13537_ : _13536_;
  assign _13539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [12] : \MSYNC_1r1w.synth.nz.mem[196] [12];
  assign _13540_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [12] : \MSYNC_1r1w.synth.nz.mem[198] [12];
  assign _13541_ = \bapg_rd.w_ptr_r [1] ? _13540_ : _13539_;
  assign _13542_ = \bapg_rd.w_ptr_r [2] ? _13541_ : _13538_;
  assign _13543_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [12] : \MSYNC_1r1w.synth.nz.mem[200] [12];
  assign _13544_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [12] : \MSYNC_1r1w.synth.nz.mem[202] [12];
  assign _13545_ = \bapg_rd.w_ptr_r [1] ? _13544_ : _13543_;
  assign _13546_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [12] : \MSYNC_1r1w.synth.nz.mem[204] [12];
  assign _13547_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [12] : \MSYNC_1r1w.synth.nz.mem[206] [12];
  assign _13548_ = \bapg_rd.w_ptr_r [1] ? _13547_ : _13546_;
  assign _13549_ = \bapg_rd.w_ptr_r [2] ? _13548_ : _13545_;
  assign _13550_ = \bapg_rd.w_ptr_r [3] ? _13549_ : _13542_;
  assign _13551_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [12] : \MSYNC_1r1w.synth.nz.mem[208] [12];
  assign _13552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [12] : \MSYNC_1r1w.synth.nz.mem[210] [12];
  assign _13553_ = \bapg_rd.w_ptr_r [1] ? _13552_ : _13551_;
  assign _13554_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [12] : \MSYNC_1r1w.synth.nz.mem[212] [12];
  assign _13555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [12] : \MSYNC_1r1w.synth.nz.mem[214] [12];
  assign _13556_ = \bapg_rd.w_ptr_r [1] ? _13555_ : _13554_;
  assign _13557_ = \bapg_rd.w_ptr_r [2] ? _13556_ : _13553_;
  assign _13558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [12] : \MSYNC_1r1w.synth.nz.mem[216] [12];
  assign _13559_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [12] : \MSYNC_1r1w.synth.nz.mem[218] [12];
  assign _13560_ = \bapg_rd.w_ptr_r [1] ? _13559_ : _13558_;
  assign _13561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [12] : \MSYNC_1r1w.synth.nz.mem[220] [12];
  assign _13562_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [12] : \MSYNC_1r1w.synth.nz.mem[222] [12];
  assign _13563_ = \bapg_rd.w_ptr_r [1] ? _13562_ : _13561_;
  assign _13564_ = \bapg_rd.w_ptr_r [2] ? _13563_ : _13560_;
  assign _13565_ = \bapg_rd.w_ptr_r [3] ? _13564_ : _13557_;
  assign _13566_ = \bapg_rd.w_ptr_r [4] ? _13565_ : _13550_;
  assign _13567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [12] : \MSYNC_1r1w.synth.nz.mem[224] [12];
  assign _13568_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [12] : \MSYNC_1r1w.synth.nz.mem[226] [12];
  assign _13569_ = \bapg_rd.w_ptr_r [1] ? _13568_ : _13567_;
  assign _13570_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [12] : \MSYNC_1r1w.synth.nz.mem[228] [12];
  assign _13571_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [12] : \MSYNC_1r1w.synth.nz.mem[230] [12];
  assign _13572_ = \bapg_rd.w_ptr_r [1] ? _13571_ : _13570_;
  assign _13573_ = \bapg_rd.w_ptr_r [2] ? _13572_ : _13569_;
  assign _13574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [12] : \MSYNC_1r1w.synth.nz.mem[232] [12];
  assign _13575_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [12] : \MSYNC_1r1w.synth.nz.mem[234] [12];
  assign _13576_ = \bapg_rd.w_ptr_r [1] ? _13575_ : _13574_;
  assign _13577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [12] : \MSYNC_1r1w.synth.nz.mem[236] [12];
  assign _13578_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [12] : \MSYNC_1r1w.synth.nz.mem[238] [12];
  assign _13579_ = \bapg_rd.w_ptr_r [1] ? _13578_ : _13577_;
  assign _13580_ = \bapg_rd.w_ptr_r [2] ? _13579_ : _13576_;
  assign _13581_ = \bapg_rd.w_ptr_r [3] ? _13580_ : _13573_;
  assign _13582_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [12] : \MSYNC_1r1w.synth.nz.mem[240] [12];
  assign _13583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [12] : \MSYNC_1r1w.synth.nz.mem[242] [12];
  assign _13584_ = \bapg_rd.w_ptr_r [1] ? _13583_ : _13582_;
  assign _13585_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [12] : \MSYNC_1r1w.synth.nz.mem[244] [12];
  assign _13586_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [12] : \MSYNC_1r1w.synth.nz.mem[246] [12];
  assign _13587_ = \bapg_rd.w_ptr_r [1] ? _13586_ : _13585_;
  assign _13588_ = \bapg_rd.w_ptr_r [2] ? _13587_ : _13584_;
  assign _13589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [12] : \MSYNC_1r1w.synth.nz.mem[248] [12];
  assign _13590_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [12] : \MSYNC_1r1w.synth.nz.mem[250] [12];
  assign _13591_ = \bapg_rd.w_ptr_r [1] ? _13590_ : _13589_;
  assign _13592_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [12] : \MSYNC_1r1w.synth.nz.mem[252] [12];
  assign _13593_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [12] : \MSYNC_1r1w.synth.nz.mem[254] [12];
  assign _13594_ = \bapg_rd.w_ptr_r [1] ? _13593_ : _13592_;
  assign _13595_ = \bapg_rd.w_ptr_r [2] ? _13594_ : _13591_;
  assign _13596_ = \bapg_rd.w_ptr_r [3] ? _13595_ : _13588_;
  assign _13597_ = \bapg_rd.w_ptr_r [4] ? _13596_ : _13581_;
  assign _13598_ = \bapg_rd.w_ptr_r [5] ? _13597_ : _13566_;
  assign _13599_ = \bapg_rd.w_ptr_r [6] ? _13598_ : _13535_;
  assign _13600_ = \bapg_rd.w_ptr_r [7] ? _13599_ : _13472_;
  assign _13601_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [12] : \MSYNC_1r1w.synth.nz.mem[256] [12];
  assign _13602_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [12] : \MSYNC_1r1w.synth.nz.mem[258] [12];
  assign _13603_ = \bapg_rd.w_ptr_r [1] ? _13602_ : _13601_;
  assign _13604_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [12] : \MSYNC_1r1w.synth.nz.mem[260] [12];
  assign _13605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [12] : \MSYNC_1r1w.synth.nz.mem[262] [12];
  assign _13606_ = \bapg_rd.w_ptr_r [1] ? _13605_ : _13604_;
  assign _13607_ = \bapg_rd.w_ptr_r [2] ? _13606_ : _13603_;
  assign _13608_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [12] : \MSYNC_1r1w.synth.nz.mem[264] [12];
  assign _13609_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [12] : \MSYNC_1r1w.synth.nz.mem[266] [12];
  assign _13610_ = \bapg_rd.w_ptr_r [1] ? _13609_ : _13608_;
  assign _13611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [12] : \MSYNC_1r1w.synth.nz.mem[268] [12];
  assign _13612_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [12] : \MSYNC_1r1w.synth.nz.mem[270] [12];
  assign _13613_ = \bapg_rd.w_ptr_r [1] ? _13612_ : _13611_;
  assign _13614_ = \bapg_rd.w_ptr_r [2] ? _13613_ : _13610_;
  assign _13615_ = \bapg_rd.w_ptr_r [3] ? _13614_ : _13607_;
  assign _13616_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [12] : \MSYNC_1r1w.synth.nz.mem[272] [12];
  assign _13617_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [12] : \MSYNC_1r1w.synth.nz.mem[274] [12];
  assign _13618_ = \bapg_rd.w_ptr_r [1] ? _13617_ : _13616_;
  assign _13619_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [12] : \MSYNC_1r1w.synth.nz.mem[276] [12];
  assign _13620_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [12] : \MSYNC_1r1w.synth.nz.mem[278] [12];
  assign _13621_ = \bapg_rd.w_ptr_r [1] ? _13620_ : _13619_;
  assign _13622_ = \bapg_rd.w_ptr_r [2] ? _13621_ : _13618_;
  assign _13623_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [12] : \MSYNC_1r1w.synth.nz.mem[280] [12];
  assign _13624_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [12] : \MSYNC_1r1w.synth.nz.mem[282] [12];
  assign _13625_ = \bapg_rd.w_ptr_r [1] ? _13624_ : _13623_;
  assign _13626_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [12] : \MSYNC_1r1w.synth.nz.mem[284] [12];
  assign _13627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [12] : \MSYNC_1r1w.synth.nz.mem[286] [12];
  assign _13628_ = \bapg_rd.w_ptr_r [1] ? _13627_ : _13626_;
  assign _13629_ = \bapg_rd.w_ptr_r [2] ? _13628_ : _13625_;
  assign _13630_ = \bapg_rd.w_ptr_r [3] ? _13629_ : _13622_;
  assign _13631_ = \bapg_rd.w_ptr_r [4] ? _13630_ : _13615_;
  assign _13632_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [12] : \MSYNC_1r1w.synth.nz.mem[288] [12];
  assign _13633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [12] : \MSYNC_1r1w.synth.nz.mem[290] [12];
  assign _13634_ = \bapg_rd.w_ptr_r [1] ? _13633_ : _13632_;
  assign _13635_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [12] : \MSYNC_1r1w.synth.nz.mem[292] [12];
  assign _13636_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [12] : \MSYNC_1r1w.synth.nz.mem[294] [12];
  assign _13637_ = \bapg_rd.w_ptr_r [1] ? _13636_ : _13635_;
  assign _13638_ = \bapg_rd.w_ptr_r [2] ? _13637_ : _13634_;
  assign _13639_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [12] : \MSYNC_1r1w.synth.nz.mem[296] [12];
  assign _13640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [12] : \MSYNC_1r1w.synth.nz.mem[298] [12];
  assign _13641_ = \bapg_rd.w_ptr_r [1] ? _13640_ : _13639_;
  assign _13642_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [12] : \MSYNC_1r1w.synth.nz.mem[300] [12];
  assign _13643_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [12] : \MSYNC_1r1w.synth.nz.mem[302] [12];
  assign _13644_ = \bapg_rd.w_ptr_r [1] ? _13643_ : _13642_;
  assign _13645_ = \bapg_rd.w_ptr_r [2] ? _13644_ : _13641_;
  assign _13646_ = \bapg_rd.w_ptr_r [3] ? _13645_ : _13638_;
  assign _13647_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [12] : \MSYNC_1r1w.synth.nz.mem[304] [12];
  assign _13648_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [12] : \MSYNC_1r1w.synth.nz.mem[306] [12];
  assign _13649_ = \bapg_rd.w_ptr_r [1] ? _13648_ : _13647_;
  assign _13650_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [12] : \MSYNC_1r1w.synth.nz.mem[308] [12];
  assign _13651_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [12] : \MSYNC_1r1w.synth.nz.mem[310] [12];
  assign _13652_ = \bapg_rd.w_ptr_r [1] ? _13651_ : _13650_;
  assign _13653_ = \bapg_rd.w_ptr_r [2] ? _13652_ : _13649_;
  assign _13654_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [12] : \MSYNC_1r1w.synth.nz.mem[312] [12];
  assign _13655_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [12] : \MSYNC_1r1w.synth.nz.mem[314] [12];
  assign _13656_ = \bapg_rd.w_ptr_r [1] ? _13655_ : _13654_;
  assign _13657_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [12] : \MSYNC_1r1w.synth.nz.mem[316] [12];
  assign _13658_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [12] : \MSYNC_1r1w.synth.nz.mem[318] [12];
  assign _13659_ = \bapg_rd.w_ptr_r [1] ? _13658_ : _13657_;
  assign _13660_ = \bapg_rd.w_ptr_r [2] ? _13659_ : _13656_;
  assign _13661_ = \bapg_rd.w_ptr_r [3] ? _13660_ : _13653_;
  assign _13662_ = \bapg_rd.w_ptr_r [4] ? _13661_ : _13646_;
  assign _13663_ = \bapg_rd.w_ptr_r [5] ? _13662_ : _13631_;
  assign _13664_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [12] : \MSYNC_1r1w.synth.nz.mem[320] [12];
  assign _13665_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [12] : \MSYNC_1r1w.synth.nz.mem[322] [12];
  assign _13666_ = \bapg_rd.w_ptr_r [1] ? _13665_ : _13664_;
  assign _13667_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [12] : \MSYNC_1r1w.synth.nz.mem[324] [12];
  assign _13668_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [12] : \MSYNC_1r1w.synth.nz.mem[326] [12];
  assign _13669_ = \bapg_rd.w_ptr_r [1] ? _13668_ : _13667_;
  assign _13670_ = \bapg_rd.w_ptr_r [2] ? _13669_ : _13666_;
  assign _13671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [12] : \MSYNC_1r1w.synth.nz.mem[328] [12];
  assign _13672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [12] : \MSYNC_1r1w.synth.nz.mem[330] [12];
  assign _13673_ = \bapg_rd.w_ptr_r [1] ? _13672_ : _13671_;
  assign _13674_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [12] : \MSYNC_1r1w.synth.nz.mem[332] [12];
  assign _13675_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [12] : \MSYNC_1r1w.synth.nz.mem[334] [12];
  assign _13676_ = \bapg_rd.w_ptr_r [1] ? _13675_ : _13674_;
  assign _13677_ = \bapg_rd.w_ptr_r [2] ? _13676_ : _13673_;
  assign _13678_ = \bapg_rd.w_ptr_r [3] ? _13677_ : _13670_;
  assign _13679_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [12] : \MSYNC_1r1w.synth.nz.mem[336] [12];
  assign _13680_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [12] : \MSYNC_1r1w.synth.nz.mem[338] [12];
  assign _13681_ = \bapg_rd.w_ptr_r [1] ? _13680_ : _13679_;
  assign _13682_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [12] : \MSYNC_1r1w.synth.nz.mem[340] [12];
  assign _13683_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [12] : \MSYNC_1r1w.synth.nz.mem[342] [12];
  assign _13684_ = \bapg_rd.w_ptr_r [1] ? _13683_ : _13682_;
  assign _13685_ = \bapg_rd.w_ptr_r [2] ? _13684_ : _13681_;
  assign _13686_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [12] : \MSYNC_1r1w.synth.nz.mem[344] [12];
  assign _13687_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [12] : \MSYNC_1r1w.synth.nz.mem[346] [12];
  assign _13688_ = \bapg_rd.w_ptr_r [1] ? _13687_ : _13686_;
  assign _13689_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [12] : \MSYNC_1r1w.synth.nz.mem[348] [12];
  assign _13690_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [12] : \MSYNC_1r1w.synth.nz.mem[350] [12];
  assign _13691_ = \bapg_rd.w_ptr_r [1] ? _13690_ : _13689_;
  assign _13692_ = \bapg_rd.w_ptr_r [2] ? _13691_ : _13688_;
  assign _13693_ = \bapg_rd.w_ptr_r [3] ? _13692_ : _13685_;
  assign _13694_ = \bapg_rd.w_ptr_r [4] ? _13693_ : _13678_;
  assign _13695_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [12] : \MSYNC_1r1w.synth.nz.mem[352] [12];
  assign _13696_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [12] : \MSYNC_1r1w.synth.nz.mem[354] [12];
  assign _13697_ = \bapg_rd.w_ptr_r [1] ? _13696_ : _13695_;
  assign _13698_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [12] : \MSYNC_1r1w.synth.nz.mem[356] [12];
  assign _13699_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [12] : \MSYNC_1r1w.synth.nz.mem[358] [12];
  assign _13700_ = \bapg_rd.w_ptr_r [1] ? _13699_ : _13698_;
  assign _13701_ = \bapg_rd.w_ptr_r [2] ? _13700_ : _13697_;
  assign _13702_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [12] : \MSYNC_1r1w.synth.nz.mem[360] [12];
  assign _13703_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [12] : \MSYNC_1r1w.synth.nz.mem[362] [12];
  assign _13704_ = \bapg_rd.w_ptr_r [1] ? _13703_ : _13702_;
  assign _13705_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [12] : \MSYNC_1r1w.synth.nz.mem[364] [12];
  assign _13706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [12] : \MSYNC_1r1w.synth.nz.mem[366] [12];
  assign _13707_ = \bapg_rd.w_ptr_r [1] ? _13706_ : _13705_;
  assign _13708_ = \bapg_rd.w_ptr_r [2] ? _13707_ : _13704_;
  assign _13709_ = \bapg_rd.w_ptr_r [3] ? _13708_ : _13701_;
  assign _13710_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [12] : \MSYNC_1r1w.synth.nz.mem[368] [12];
  assign _13711_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [12] : \MSYNC_1r1w.synth.nz.mem[370] [12];
  assign _13712_ = \bapg_rd.w_ptr_r [1] ? _13711_ : _13710_;
  assign _13713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [12] : \MSYNC_1r1w.synth.nz.mem[372] [12];
  assign _13714_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [12] : \MSYNC_1r1w.synth.nz.mem[374] [12];
  assign _13715_ = \bapg_rd.w_ptr_r [1] ? _13714_ : _13713_;
  assign _13716_ = \bapg_rd.w_ptr_r [2] ? _13715_ : _13712_;
  assign _13717_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [12] : \MSYNC_1r1w.synth.nz.mem[376] [12];
  assign _13718_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [12] : \MSYNC_1r1w.synth.nz.mem[378] [12];
  assign _13719_ = \bapg_rd.w_ptr_r [1] ? _13718_ : _13717_;
  assign _13720_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [12] : \MSYNC_1r1w.synth.nz.mem[380] [12];
  assign _13721_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [12] : \MSYNC_1r1w.synth.nz.mem[382] [12];
  assign _13722_ = \bapg_rd.w_ptr_r [1] ? _13721_ : _13720_;
  assign _13723_ = \bapg_rd.w_ptr_r [2] ? _13722_ : _13719_;
  assign _13724_ = \bapg_rd.w_ptr_r [3] ? _13723_ : _13716_;
  assign _13725_ = \bapg_rd.w_ptr_r [4] ? _13724_ : _13709_;
  assign _13726_ = \bapg_rd.w_ptr_r [5] ? _13725_ : _13694_;
  assign _13727_ = \bapg_rd.w_ptr_r [6] ? _13726_ : _13663_;
  assign _13728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [12] : \MSYNC_1r1w.synth.nz.mem[384] [12];
  assign _13729_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [12] : \MSYNC_1r1w.synth.nz.mem[386] [12];
  assign _13730_ = \bapg_rd.w_ptr_r [1] ? _13729_ : _13728_;
  assign _13731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [12] : \MSYNC_1r1w.synth.nz.mem[388] [12];
  assign _13732_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [12] : \MSYNC_1r1w.synth.nz.mem[390] [12];
  assign _13733_ = \bapg_rd.w_ptr_r [1] ? _13732_ : _13731_;
  assign _13734_ = \bapg_rd.w_ptr_r [2] ? _13733_ : _13730_;
  assign _13735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [12] : \MSYNC_1r1w.synth.nz.mem[392] [12];
  assign _13736_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [12] : \MSYNC_1r1w.synth.nz.mem[394] [12];
  assign _13737_ = \bapg_rd.w_ptr_r [1] ? _13736_ : _13735_;
  assign _13738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [12] : \MSYNC_1r1w.synth.nz.mem[396] [12];
  assign _13739_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [12] : \MSYNC_1r1w.synth.nz.mem[398] [12];
  assign _13740_ = \bapg_rd.w_ptr_r [1] ? _13739_ : _13738_;
  assign _13741_ = \bapg_rd.w_ptr_r [2] ? _13740_ : _13737_;
  assign _13742_ = \bapg_rd.w_ptr_r [3] ? _13741_ : _13734_;
  assign _13743_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [12] : \MSYNC_1r1w.synth.nz.mem[400] [12];
  assign _13744_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [12] : \MSYNC_1r1w.synth.nz.mem[402] [12];
  assign _13745_ = \bapg_rd.w_ptr_r [1] ? _13744_ : _13743_;
  assign _13746_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [12] : \MSYNC_1r1w.synth.nz.mem[404] [12];
  assign _13747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [12] : \MSYNC_1r1w.synth.nz.mem[406] [12];
  assign _13748_ = \bapg_rd.w_ptr_r [1] ? _13747_ : _13746_;
  assign _13749_ = \bapg_rd.w_ptr_r [2] ? _13748_ : _13745_;
  assign _13750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [12] : \MSYNC_1r1w.synth.nz.mem[408] [12];
  assign _13751_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [12] : \MSYNC_1r1w.synth.nz.mem[410] [12];
  assign _13752_ = \bapg_rd.w_ptr_r [1] ? _13751_ : _13750_;
  assign _13753_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [12] : \MSYNC_1r1w.synth.nz.mem[412] [12];
  assign _13754_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [12] : \MSYNC_1r1w.synth.nz.mem[414] [12];
  assign _13755_ = \bapg_rd.w_ptr_r [1] ? _13754_ : _13753_;
  assign _13756_ = \bapg_rd.w_ptr_r [2] ? _13755_ : _13752_;
  assign _13757_ = \bapg_rd.w_ptr_r [3] ? _13756_ : _13749_;
  assign _13758_ = \bapg_rd.w_ptr_r [4] ? _13757_ : _13742_;
  assign _13759_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [12] : \MSYNC_1r1w.synth.nz.mem[416] [12];
  assign _13760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [12] : \MSYNC_1r1w.synth.nz.mem[418] [12];
  assign _13761_ = \bapg_rd.w_ptr_r [1] ? _13760_ : _13759_;
  assign _13762_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [12] : \MSYNC_1r1w.synth.nz.mem[420] [12];
  assign _13763_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [12] : \MSYNC_1r1w.synth.nz.mem[422] [12];
  assign _13764_ = \bapg_rd.w_ptr_r [1] ? _13763_ : _13762_;
  assign _13765_ = \bapg_rd.w_ptr_r [2] ? _13764_ : _13761_;
  assign _13766_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [12] : \MSYNC_1r1w.synth.nz.mem[424] [12];
  assign _13767_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [12] : \MSYNC_1r1w.synth.nz.mem[426] [12];
  assign _13768_ = \bapg_rd.w_ptr_r [1] ? _13767_ : _13766_;
  assign _13769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [12] : \MSYNC_1r1w.synth.nz.mem[428] [12];
  assign _13770_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [12] : \MSYNC_1r1w.synth.nz.mem[430] [12];
  assign _13771_ = \bapg_rd.w_ptr_r [1] ? _13770_ : _13769_;
  assign _13772_ = \bapg_rd.w_ptr_r [2] ? _13771_ : _13768_;
  assign _13773_ = \bapg_rd.w_ptr_r [3] ? _13772_ : _13765_;
  assign _13774_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [12] : \MSYNC_1r1w.synth.nz.mem[432] [12];
  assign _13775_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [12] : \MSYNC_1r1w.synth.nz.mem[434] [12];
  assign _13776_ = \bapg_rd.w_ptr_r [1] ? _13775_ : _13774_;
  assign _13777_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [12] : \MSYNC_1r1w.synth.nz.mem[436] [12];
  assign _13778_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [12] : \MSYNC_1r1w.synth.nz.mem[438] [12];
  assign _13779_ = \bapg_rd.w_ptr_r [1] ? _13778_ : _13777_;
  assign _13780_ = \bapg_rd.w_ptr_r [2] ? _13779_ : _13776_;
  assign _13781_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [12] : \MSYNC_1r1w.synth.nz.mem[440] [12];
  assign _13782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [12] : \MSYNC_1r1w.synth.nz.mem[442] [12];
  assign _13783_ = \bapg_rd.w_ptr_r [1] ? _13782_ : _13781_;
  assign _13784_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [12] : \MSYNC_1r1w.synth.nz.mem[444] [12];
  assign _13785_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [12] : \MSYNC_1r1w.synth.nz.mem[446] [12];
  assign _13786_ = \bapg_rd.w_ptr_r [1] ? _13785_ : _13784_;
  assign _13787_ = \bapg_rd.w_ptr_r [2] ? _13786_ : _13783_;
  assign _13788_ = \bapg_rd.w_ptr_r [3] ? _13787_ : _13780_;
  assign _13789_ = \bapg_rd.w_ptr_r [4] ? _13788_ : _13773_;
  assign _13790_ = \bapg_rd.w_ptr_r [5] ? _13789_ : _13758_;
  assign _13791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [12] : \MSYNC_1r1w.synth.nz.mem[448] [12];
  assign _13792_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [12] : \MSYNC_1r1w.synth.nz.mem[450] [12];
  assign _13793_ = \bapg_rd.w_ptr_r [1] ? _13792_ : _13791_;
  assign _13794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [12] : \MSYNC_1r1w.synth.nz.mem[452] [12];
  assign _13795_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [12] : \MSYNC_1r1w.synth.nz.mem[454] [12];
  assign _13796_ = \bapg_rd.w_ptr_r [1] ? _13795_ : _13794_;
  assign _13797_ = \bapg_rd.w_ptr_r [2] ? _13796_ : _13793_;
  assign _13798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [12] : \MSYNC_1r1w.synth.nz.mem[456] [12];
  assign _13799_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [12] : \MSYNC_1r1w.synth.nz.mem[458] [12];
  assign _13800_ = \bapg_rd.w_ptr_r [1] ? _13799_ : _13798_;
  assign _13801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [12] : \MSYNC_1r1w.synth.nz.mem[460] [12];
  assign _13802_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [12] : \MSYNC_1r1w.synth.nz.mem[462] [12];
  assign _13803_ = \bapg_rd.w_ptr_r [1] ? _13802_ : _13801_;
  assign _13804_ = \bapg_rd.w_ptr_r [2] ? _13803_ : _13800_;
  assign _13805_ = \bapg_rd.w_ptr_r [3] ? _13804_ : _13797_;
  assign _13806_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [12] : \MSYNC_1r1w.synth.nz.mem[464] [12];
  assign _13807_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [12] : \MSYNC_1r1w.synth.nz.mem[466] [12];
  assign _13808_ = \bapg_rd.w_ptr_r [1] ? _13807_ : _13806_;
  assign _13809_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [12] : \MSYNC_1r1w.synth.nz.mem[468] [12];
  assign _13810_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [12] : \MSYNC_1r1w.synth.nz.mem[470] [12];
  assign _13811_ = \bapg_rd.w_ptr_r [1] ? _13810_ : _13809_;
  assign _13812_ = \bapg_rd.w_ptr_r [2] ? _13811_ : _13808_;
  assign _13813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [12] : \MSYNC_1r1w.synth.nz.mem[472] [12];
  assign _13814_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [12] : \MSYNC_1r1w.synth.nz.mem[474] [12];
  assign _13815_ = \bapg_rd.w_ptr_r [1] ? _13814_ : _13813_;
  assign _13816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [12] : \MSYNC_1r1w.synth.nz.mem[476] [12];
  assign _13817_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [12] : \MSYNC_1r1w.synth.nz.mem[478] [12];
  assign _13818_ = \bapg_rd.w_ptr_r [1] ? _13817_ : _13816_;
  assign _13819_ = \bapg_rd.w_ptr_r [2] ? _13818_ : _13815_;
  assign _13820_ = \bapg_rd.w_ptr_r [3] ? _13819_ : _13812_;
  assign _13821_ = \bapg_rd.w_ptr_r [4] ? _13820_ : _13805_;
  assign _13822_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [12] : \MSYNC_1r1w.synth.nz.mem[480] [12];
  assign _13823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [12] : \MSYNC_1r1w.synth.nz.mem[482] [12];
  assign _13824_ = \bapg_rd.w_ptr_r [1] ? _13823_ : _13822_;
  assign _13825_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [12] : \MSYNC_1r1w.synth.nz.mem[484] [12];
  assign _13826_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [12] : \MSYNC_1r1w.synth.nz.mem[486] [12];
  assign _13827_ = \bapg_rd.w_ptr_r [1] ? _13826_ : _13825_;
  assign _13828_ = \bapg_rd.w_ptr_r [2] ? _13827_ : _13824_;
  assign _13829_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [12] : \MSYNC_1r1w.synth.nz.mem[488] [12];
  assign _13830_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [12] : \MSYNC_1r1w.synth.nz.mem[490] [12];
  assign _13831_ = \bapg_rd.w_ptr_r [1] ? _13830_ : _13829_;
  assign _13832_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [12] : \MSYNC_1r1w.synth.nz.mem[492] [12];
  assign _13833_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [12] : \MSYNC_1r1w.synth.nz.mem[494] [12];
  assign _13834_ = \bapg_rd.w_ptr_r [1] ? _13833_ : _13832_;
  assign _13835_ = \bapg_rd.w_ptr_r [2] ? _13834_ : _13831_;
  assign _13836_ = \bapg_rd.w_ptr_r [3] ? _13835_ : _13828_;
  assign _13837_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [12] : \MSYNC_1r1w.synth.nz.mem[496] [12];
  assign _13838_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [12] : \MSYNC_1r1w.synth.nz.mem[498] [12];
  assign _13839_ = \bapg_rd.w_ptr_r [1] ? _13838_ : _13837_;
  assign _13840_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [12] : \MSYNC_1r1w.synth.nz.mem[500] [12];
  assign _13841_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [12] : \MSYNC_1r1w.synth.nz.mem[502] [12];
  assign _13842_ = \bapg_rd.w_ptr_r [1] ? _13841_ : _13840_;
  assign _13843_ = \bapg_rd.w_ptr_r [2] ? _13842_ : _13839_;
  assign _13844_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [12] : \MSYNC_1r1w.synth.nz.mem[504] [12];
  assign _13845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [12] : \MSYNC_1r1w.synth.nz.mem[506] [12];
  assign _13846_ = \bapg_rd.w_ptr_r [1] ? _13845_ : _13844_;
  assign _13847_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [12] : \MSYNC_1r1w.synth.nz.mem[508] [12];
  assign _13848_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [12] : \MSYNC_1r1w.synth.nz.mem[510] [12];
  assign _13849_ = \bapg_rd.w_ptr_r [1] ? _13848_ : _13847_;
  assign _13850_ = \bapg_rd.w_ptr_r [2] ? _13849_ : _13846_;
  assign _13851_ = \bapg_rd.w_ptr_r [3] ? _13850_ : _13843_;
  assign _13852_ = \bapg_rd.w_ptr_r [4] ? _13851_ : _13836_;
  assign _13853_ = \bapg_rd.w_ptr_r [5] ? _13852_ : _13821_;
  assign _13854_ = \bapg_rd.w_ptr_r [6] ? _13853_ : _13790_;
  assign _13855_ = \bapg_rd.w_ptr_r [7] ? _13854_ : _13727_;
  assign _13856_ = \bapg_rd.w_ptr_r [8] ? _13855_ : _13600_;
  assign _13857_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [12] : \MSYNC_1r1w.synth.nz.mem[512] [12];
  assign _13858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [12] : \MSYNC_1r1w.synth.nz.mem[514] [12];
  assign _13859_ = \bapg_rd.w_ptr_r [1] ? _13858_ : _13857_;
  assign _13860_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [12] : \MSYNC_1r1w.synth.nz.mem[516] [12];
  assign _13861_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [12] : \MSYNC_1r1w.synth.nz.mem[518] [12];
  assign _13862_ = \bapg_rd.w_ptr_r [1] ? _13861_ : _13860_;
  assign _13863_ = \bapg_rd.w_ptr_r [2] ? _13862_ : _13859_;
  assign _13864_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [12] : \MSYNC_1r1w.synth.nz.mem[520] [12];
  assign _13865_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [12] : \MSYNC_1r1w.synth.nz.mem[522] [12];
  assign _13866_ = \bapg_rd.w_ptr_r [1] ? _13865_ : _13864_;
  assign _13867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [12] : \MSYNC_1r1w.synth.nz.mem[524] [12];
  assign _13868_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [12] : \MSYNC_1r1w.synth.nz.mem[526] [12];
  assign _13869_ = \bapg_rd.w_ptr_r [1] ? _13868_ : _13867_;
  assign _13870_ = \bapg_rd.w_ptr_r [2] ? _13869_ : _13866_;
  assign _13871_ = \bapg_rd.w_ptr_r [3] ? _13870_ : _13863_;
  assign _13872_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [12] : \MSYNC_1r1w.synth.nz.mem[528] [12];
  assign _13873_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [12] : \MSYNC_1r1w.synth.nz.mem[530] [12];
  assign _13874_ = \bapg_rd.w_ptr_r [1] ? _13873_ : _13872_;
  assign _13875_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [12] : \MSYNC_1r1w.synth.nz.mem[532] [12];
  assign _13876_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [12] : \MSYNC_1r1w.synth.nz.mem[534] [12];
  assign _13877_ = \bapg_rd.w_ptr_r [1] ? _13876_ : _13875_;
  assign _13878_ = \bapg_rd.w_ptr_r [2] ? _13877_ : _13874_;
  assign _13879_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [12] : \MSYNC_1r1w.synth.nz.mem[536] [12];
  assign _13880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [12] : \MSYNC_1r1w.synth.nz.mem[538] [12];
  assign _13881_ = \bapg_rd.w_ptr_r [1] ? _13880_ : _13879_;
  assign _13882_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [12] : \MSYNC_1r1w.synth.nz.mem[540] [12];
  assign _13883_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [12] : \MSYNC_1r1w.synth.nz.mem[542] [12];
  assign _13884_ = \bapg_rd.w_ptr_r [1] ? _13883_ : _13882_;
  assign _13885_ = \bapg_rd.w_ptr_r [2] ? _13884_ : _13881_;
  assign _13886_ = \bapg_rd.w_ptr_r [3] ? _13885_ : _13878_;
  assign _13887_ = \bapg_rd.w_ptr_r [4] ? _13886_ : _13871_;
  assign _13888_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [12] : \MSYNC_1r1w.synth.nz.mem[544] [12];
  assign _13889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [12] : \MSYNC_1r1w.synth.nz.mem[546] [12];
  assign _13890_ = \bapg_rd.w_ptr_r [1] ? _13889_ : _13888_;
  assign _13891_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [12] : \MSYNC_1r1w.synth.nz.mem[548] [12];
  assign _13892_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [12] : \MSYNC_1r1w.synth.nz.mem[550] [12];
  assign _13893_ = \bapg_rd.w_ptr_r [1] ? _13892_ : _13891_;
  assign _13894_ = \bapg_rd.w_ptr_r [2] ? _13893_ : _13890_;
  assign _13895_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [12] : \MSYNC_1r1w.synth.nz.mem[552] [12];
  assign _13896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [12] : \MSYNC_1r1w.synth.nz.mem[554] [12];
  assign _13897_ = \bapg_rd.w_ptr_r [1] ? _13896_ : _13895_;
  assign _13898_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [12] : \MSYNC_1r1w.synth.nz.mem[556] [12];
  assign _13899_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [12] : \MSYNC_1r1w.synth.nz.mem[558] [12];
  assign _13900_ = \bapg_rd.w_ptr_r [1] ? _13899_ : _13898_;
  assign _13901_ = \bapg_rd.w_ptr_r [2] ? _13900_ : _13897_;
  assign _13902_ = \bapg_rd.w_ptr_r [3] ? _13901_ : _13894_;
  assign _13903_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [12] : \MSYNC_1r1w.synth.nz.mem[560] [12];
  assign _13904_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [12] : \MSYNC_1r1w.synth.nz.mem[562] [12];
  assign _13905_ = \bapg_rd.w_ptr_r [1] ? _13904_ : _13903_;
  assign _13906_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [12] : \MSYNC_1r1w.synth.nz.mem[564] [12];
  assign _13907_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [12] : \MSYNC_1r1w.synth.nz.mem[566] [12];
  assign _13908_ = \bapg_rd.w_ptr_r [1] ? _13907_ : _13906_;
  assign _13909_ = \bapg_rd.w_ptr_r [2] ? _13908_ : _13905_;
  assign _13910_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [12] : \MSYNC_1r1w.synth.nz.mem[568] [12];
  assign _13911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [12] : \MSYNC_1r1w.synth.nz.mem[570] [12];
  assign _13912_ = \bapg_rd.w_ptr_r [1] ? _13911_ : _13910_;
  assign _13913_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [12] : \MSYNC_1r1w.synth.nz.mem[572] [12];
  assign _13914_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [12] : \MSYNC_1r1w.synth.nz.mem[574] [12];
  assign _13915_ = \bapg_rd.w_ptr_r [1] ? _13914_ : _13913_;
  assign _13916_ = \bapg_rd.w_ptr_r [2] ? _13915_ : _13912_;
  assign _13917_ = \bapg_rd.w_ptr_r [3] ? _13916_ : _13909_;
  assign _13918_ = \bapg_rd.w_ptr_r [4] ? _13917_ : _13902_;
  assign _13919_ = \bapg_rd.w_ptr_r [5] ? _13918_ : _13887_;
  assign _13920_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [12] : \MSYNC_1r1w.synth.nz.mem[576] [12];
  assign _13921_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [12] : \MSYNC_1r1w.synth.nz.mem[578] [12];
  assign _13922_ = \bapg_rd.w_ptr_r [1] ? _13921_ : _13920_;
  assign _13923_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [12] : \MSYNC_1r1w.synth.nz.mem[580] [12];
  assign _13924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [12] : \MSYNC_1r1w.synth.nz.mem[582] [12];
  assign _13925_ = \bapg_rd.w_ptr_r [1] ? _13924_ : _13923_;
  assign _13926_ = \bapg_rd.w_ptr_r [2] ? _13925_ : _13922_;
  assign _13927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [12] : \MSYNC_1r1w.synth.nz.mem[584] [12];
  assign _13928_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [12] : \MSYNC_1r1w.synth.nz.mem[586] [12];
  assign _13929_ = \bapg_rd.w_ptr_r [1] ? _13928_ : _13927_;
  assign _13930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [12] : \MSYNC_1r1w.synth.nz.mem[588] [12];
  assign _13931_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [12] : \MSYNC_1r1w.synth.nz.mem[590] [12];
  assign _13932_ = \bapg_rd.w_ptr_r [1] ? _13931_ : _13930_;
  assign _13933_ = \bapg_rd.w_ptr_r [2] ? _13932_ : _13929_;
  assign _13934_ = \bapg_rd.w_ptr_r [3] ? _13933_ : _13926_;
  assign _13935_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [12] : \MSYNC_1r1w.synth.nz.mem[592] [12];
  assign _13936_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [12] : \MSYNC_1r1w.synth.nz.mem[594] [12];
  assign _13937_ = \bapg_rd.w_ptr_r [1] ? _13936_ : _13935_;
  assign _13938_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [12] : \MSYNC_1r1w.synth.nz.mem[596] [12];
  assign _13939_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [12] : \MSYNC_1r1w.synth.nz.mem[598] [12];
  assign _13940_ = \bapg_rd.w_ptr_r [1] ? _13939_ : _13938_;
  assign _13941_ = \bapg_rd.w_ptr_r [2] ? _13940_ : _13937_;
  assign _13942_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [12] : \MSYNC_1r1w.synth.nz.mem[600] [12];
  assign _13943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [12] : \MSYNC_1r1w.synth.nz.mem[602] [12];
  assign _13944_ = \bapg_rd.w_ptr_r [1] ? _13943_ : _13942_;
  assign _13945_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [12] : \MSYNC_1r1w.synth.nz.mem[604] [12];
  assign _13946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [12] : \MSYNC_1r1w.synth.nz.mem[606] [12];
  assign _13947_ = \bapg_rd.w_ptr_r [1] ? _13946_ : _13945_;
  assign _13948_ = \bapg_rd.w_ptr_r [2] ? _13947_ : _13944_;
  assign _13949_ = \bapg_rd.w_ptr_r [3] ? _13948_ : _13941_;
  assign _13950_ = \bapg_rd.w_ptr_r [4] ? _13949_ : _13934_;
  assign _13951_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [12] : \MSYNC_1r1w.synth.nz.mem[608] [12];
  assign _13952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [12] : \MSYNC_1r1w.synth.nz.mem[610] [12];
  assign _13953_ = \bapg_rd.w_ptr_r [1] ? _13952_ : _13951_;
  assign _13954_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [12] : \MSYNC_1r1w.synth.nz.mem[612] [12];
  assign _13955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [12] : \MSYNC_1r1w.synth.nz.mem[614] [12];
  assign _13956_ = \bapg_rd.w_ptr_r [1] ? _13955_ : _13954_;
  assign _13957_ = \bapg_rd.w_ptr_r [2] ? _13956_ : _13953_;
  assign _13958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [12] : \MSYNC_1r1w.synth.nz.mem[616] [12];
  assign _13959_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [12] : \MSYNC_1r1w.synth.nz.mem[618] [12];
  assign _13960_ = \bapg_rd.w_ptr_r [1] ? _13959_ : _13958_;
  assign _13961_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [12] : \MSYNC_1r1w.synth.nz.mem[620] [12];
  assign _13962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [12] : \MSYNC_1r1w.synth.nz.mem[622] [12];
  assign _13963_ = \bapg_rd.w_ptr_r [1] ? _13962_ : _13961_;
  assign _13964_ = \bapg_rd.w_ptr_r [2] ? _13963_ : _13960_;
  assign _13965_ = \bapg_rd.w_ptr_r [3] ? _13964_ : _13957_;
  assign _13966_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [12] : \MSYNC_1r1w.synth.nz.mem[624] [12];
  assign _13967_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [12] : \MSYNC_1r1w.synth.nz.mem[626] [12];
  assign _13968_ = \bapg_rd.w_ptr_r [1] ? _13967_ : _13966_;
  assign _13969_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [12] : \MSYNC_1r1w.synth.nz.mem[628] [12];
  assign _13970_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [12] : \MSYNC_1r1w.synth.nz.mem[630] [12];
  assign _13971_ = \bapg_rd.w_ptr_r [1] ? _13970_ : _13969_;
  assign _13972_ = \bapg_rd.w_ptr_r [2] ? _13971_ : _13968_;
  assign _13973_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [12] : \MSYNC_1r1w.synth.nz.mem[632] [12];
  assign _13974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [12] : \MSYNC_1r1w.synth.nz.mem[634] [12];
  assign _13975_ = \bapg_rd.w_ptr_r [1] ? _13974_ : _13973_;
  assign _13976_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [12] : \MSYNC_1r1w.synth.nz.mem[636] [12];
  assign _13977_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [12] : \MSYNC_1r1w.synth.nz.mem[638] [12];
  assign _13978_ = \bapg_rd.w_ptr_r [1] ? _13977_ : _13976_;
  assign _13979_ = \bapg_rd.w_ptr_r [2] ? _13978_ : _13975_;
  assign _13980_ = \bapg_rd.w_ptr_r [3] ? _13979_ : _13972_;
  assign _13981_ = \bapg_rd.w_ptr_r [4] ? _13980_ : _13965_;
  assign _13982_ = \bapg_rd.w_ptr_r [5] ? _13981_ : _13950_;
  assign _13983_ = \bapg_rd.w_ptr_r [6] ? _13982_ : _13919_;
  assign _13984_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [12] : \MSYNC_1r1w.synth.nz.mem[640] [12];
  assign _13985_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [12] : \MSYNC_1r1w.synth.nz.mem[642] [12];
  assign _13986_ = \bapg_rd.w_ptr_r [1] ? _13985_ : _13984_;
  assign _13987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [12] : \MSYNC_1r1w.synth.nz.mem[644] [12];
  assign _13988_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [12] : \MSYNC_1r1w.synth.nz.mem[646] [12];
  assign _13989_ = \bapg_rd.w_ptr_r [1] ? _13988_ : _13987_;
  assign _13990_ = \bapg_rd.w_ptr_r [2] ? _13989_ : _13986_;
  assign _13991_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [12] : \MSYNC_1r1w.synth.nz.mem[648] [12];
  assign _13992_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [12] : \MSYNC_1r1w.synth.nz.mem[650] [12];
  assign _13993_ = \bapg_rd.w_ptr_r [1] ? _13992_ : _13991_;
  assign _13994_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [12] : \MSYNC_1r1w.synth.nz.mem[652] [12];
  assign _13995_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [12] : \MSYNC_1r1w.synth.nz.mem[654] [12];
  assign _13996_ = \bapg_rd.w_ptr_r [1] ? _13995_ : _13994_;
  assign _13997_ = \bapg_rd.w_ptr_r [2] ? _13996_ : _13993_;
  assign _13998_ = \bapg_rd.w_ptr_r [3] ? _13997_ : _13990_;
  assign _13999_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [12] : \MSYNC_1r1w.synth.nz.mem[656] [12];
  assign _14000_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [12] : \MSYNC_1r1w.synth.nz.mem[658] [12];
  assign _14001_ = \bapg_rd.w_ptr_r [1] ? _14000_ : _13999_;
  assign _14002_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [12] : \MSYNC_1r1w.synth.nz.mem[660] [12];
  assign _14003_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [12] : \MSYNC_1r1w.synth.nz.mem[662] [12];
  assign _14004_ = \bapg_rd.w_ptr_r [1] ? _14003_ : _14002_;
  assign _14005_ = \bapg_rd.w_ptr_r [2] ? _14004_ : _14001_;
  assign _14006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [12] : \MSYNC_1r1w.synth.nz.mem[664] [12];
  assign _14007_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [12] : \MSYNC_1r1w.synth.nz.mem[666] [12];
  assign _14008_ = \bapg_rd.w_ptr_r [1] ? _14007_ : _14006_;
  assign _14009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [12] : \MSYNC_1r1w.synth.nz.mem[668] [12];
  assign _14010_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [12] : \MSYNC_1r1w.synth.nz.mem[670] [12];
  assign _14011_ = \bapg_rd.w_ptr_r [1] ? _14010_ : _14009_;
  assign _14012_ = \bapg_rd.w_ptr_r [2] ? _14011_ : _14008_;
  assign _14013_ = \bapg_rd.w_ptr_r [3] ? _14012_ : _14005_;
  assign _14014_ = \bapg_rd.w_ptr_r [4] ? _14013_ : _13998_;
  assign _14015_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [12] : \MSYNC_1r1w.synth.nz.mem[672] [12];
  assign _14016_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [12] : \MSYNC_1r1w.synth.nz.mem[674] [12];
  assign _14017_ = \bapg_rd.w_ptr_r [1] ? _14016_ : _14015_;
  assign _14018_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [12] : \MSYNC_1r1w.synth.nz.mem[676] [12];
  assign _14019_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [12] : \MSYNC_1r1w.synth.nz.mem[678] [12];
  assign _14020_ = \bapg_rd.w_ptr_r [1] ? _14019_ : _14018_;
  assign _14021_ = \bapg_rd.w_ptr_r [2] ? _14020_ : _14017_;
  assign _14022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [12] : \MSYNC_1r1w.synth.nz.mem[680] [12];
  assign _14023_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [12] : \MSYNC_1r1w.synth.nz.mem[682] [12];
  assign _14024_ = \bapg_rd.w_ptr_r [1] ? _14023_ : _14022_;
  assign _14025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [12] : \MSYNC_1r1w.synth.nz.mem[684] [12];
  assign _14026_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [12] : \MSYNC_1r1w.synth.nz.mem[686] [12];
  assign _14027_ = \bapg_rd.w_ptr_r [1] ? _14026_ : _14025_;
  assign _14028_ = \bapg_rd.w_ptr_r [2] ? _14027_ : _14024_;
  assign _14029_ = \bapg_rd.w_ptr_r [3] ? _14028_ : _14021_;
  assign _14030_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [12] : \MSYNC_1r1w.synth.nz.mem[688] [12];
  assign _14031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [12] : \MSYNC_1r1w.synth.nz.mem[690] [12];
  assign _14032_ = \bapg_rd.w_ptr_r [1] ? _14031_ : _14030_;
  assign _14033_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [12] : \MSYNC_1r1w.synth.nz.mem[692] [12];
  assign _14034_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [12] : \MSYNC_1r1w.synth.nz.mem[694] [12];
  assign _14035_ = \bapg_rd.w_ptr_r [1] ? _14034_ : _14033_;
  assign _14036_ = \bapg_rd.w_ptr_r [2] ? _14035_ : _14032_;
  assign _14037_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [12] : \MSYNC_1r1w.synth.nz.mem[696] [12];
  assign _14038_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [12] : \MSYNC_1r1w.synth.nz.mem[698] [12];
  assign _14039_ = \bapg_rd.w_ptr_r [1] ? _14038_ : _14037_;
  assign _14040_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [12] : \MSYNC_1r1w.synth.nz.mem[700] [12];
  assign _14041_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [12] : \MSYNC_1r1w.synth.nz.mem[702] [12];
  assign _14042_ = \bapg_rd.w_ptr_r [1] ? _14041_ : _14040_;
  assign _14043_ = \bapg_rd.w_ptr_r [2] ? _14042_ : _14039_;
  assign _14044_ = \bapg_rd.w_ptr_r [3] ? _14043_ : _14036_;
  assign _14045_ = \bapg_rd.w_ptr_r [4] ? _14044_ : _14029_;
  assign _14046_ = \bapg_rd.w_ptr_r [5] ? _14045_ : _14014_;
  assign _14047_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [12] : \MSYNC_1r1w.synth.nz.mem[704] [12];
  assign _14048_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [12] : \MSYNC_1r1w.synth.nz.mem[706] [12];
  assign _14049_ = \bapg_rd.w_ptr_r [1] ? _14048_ : _14047_;
  assign _14050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [12] : \MSYNC_1r1w.synth.nz.mem[708] [12];
  assign _14051_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [12] : \MSYNC_1r1w.synth.nz.mem[710] [12];
  assign _14052_ = \bapg_rd.w_ptr_r [1] ? _14051_ : _14050_;
  assign _14053_ = \bapg_rd.w_ptr_r [2] ? _14052_ : _14049_;
  assign _14054_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [12] : \MSYNC_1r1w.synth.nz.mem[712] [12];
  assign _14055_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [12] : \MSYNC_1r1w.synth.nz.mem[714] [12];
  assign _14056_ = \bapg_rd.w_ptr_r [1] ? _14055_ : _14054_;
  assign _14057_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [12] : \MSYNC_1r1w.synth.nz.mem[716] [12];
  assign _14058_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [12] : \MSYNC_1r1w.synth.nz.mem[718] [12];
  assign _14059_ = \bapg_rd.w_ptr_r [1] ? _14058_ : _14057_;
  assign _14060_ = \bapg_rd.w_ptr_r [2] ? _14059_ : _14056_;
  assign _14061_ = \bapg_rd.w_ptr_r [3] ? _14060_ : _14053_;
  assign _14062_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [12] : \MSYNC_1r1w.synth.nz.mem[720] [12];
  assign _14063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [12] : \MSYNC_1r1w.synth.nz.mem[722] [12];
  assign _14064_ = \bapg_rd.w_ptr_r [1] ? _14063_ : _14062_;
  assign _14065_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [12] : \MSYNC_1r1w.synth.nz.mem[724] [12];
  assign _14066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [12] : \MSYNC_1r1w.synth.nz.mem[726] [12];
  assign _14067_ = \bapg_rd.w_ptr_r [1] ? _14066_ : _14065_;
  assign _14068_ = \bapg_rd.w_ptr_r [2] ? _14067_ : _14064_;
  assign _14069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [12] : \MSYNC_1r1w.synth.nz.mem[728] [12];
  assign _14070_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [12] : \MSYNC_1r1w.synth.nz.mem[730] [12];
  assign _14071_ = \bapg_rd.w_ptr_r [1] ? _14070_ : _14069_;
  assign _14072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [12] : \MSYNC_1r1w.synth.nz.mem[732] [12];
  assign _14073_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [12] : \MSYNC_1r1w.synth.nz.mem[734] [12];
  assign _14074_ = \bapg_rd.w_ptr_r [1] ? _14073_ : _14072_;
  assign _14075_ = \bapg_rd.w_ptr_r [2] ? _14074_ : _14071_;
  assign _14076_ = \bapg_rd.w_ptr_r [3] ? _14075_ : _14068_;
  assign _14077_ = \bapg_rd.w_ptr_r [4] ? _14076_ : _14061_;
  assign _14078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [12] : \MSYNC_1r1w.synth.nz.mem[736] [12];
  assign _14079_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [12] : \MSYNC_1r1w.synth.nz.mem[738] [12];
  assign _14080_ = \bapg_rd.w_ptr_r [1] ? _14079_ : _14078_;
  assign _14081_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [12] : \MSYNC_1r1w.synth.nz.mem[740] [12];
  assign _14082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [12] : \MSYNC_1r1w.synth.nz.mem[742] [12];
  assign _14083_ = \bapg_rd.w_ptr_r [1] ? _14082_ : _14081_;
  assign _14084_ = \bapg_rd.w_ptr_r [2] ? _14083_ : _14080_;
  assign _14085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [12] : \MSYNC_1r1w.synth.nz.mem[744] [12];
  assign _14086_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [12] : \MSYNC_1r1w.synth.nz.mem[746] [12];
  assign _14087_ = \bapg_rd.w_ptr_r [1] ? _14086_ : _14085_;
  assign _14088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [12] : \MSYNC_1r1w.synth.nz.mem[748] [12];
  assign _14089_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [12] : \MSYNC_1r1w.synth.nz.mem[750] [12];
  assign _14090_ = \bapg_rd.w_ptr_r [1] ? _14089_ : _14088_;
  assign _14091_ = \bapg_rd.w_ptr_r [2] ? _14090_ : _14087_;
  assign _14092_ = \bapg_rd.w_ptr_r [3] ? _14091_ : _14084_;
  assign _14093_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [12] : \MSYNC_1r1w.synth.nz.mem[752] [12];
  assign _14094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [12] : \MSYNC_1r1w.synth.nz.mem[754] [12];
  assign _14095_ = \bapg_rd.w_ptr_r [1] ? _14094_ : _14093_;
  assign _14096_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [12] : \MSYNC_1r1w.synth.nz.mem[756] [12];
  assign _14097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [12] : \MSYNC_1r1w.synth.nz.mem[758] [12];
  assign _14098_ = \bapg_rd.w_ptr_r [1] ? _14097_ : _14096_;
  assign _14099_ = \bapg_rd.w_ptr_r [2] ? _14098_ : _14095_;
  assign _14100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [12] : \MSYNC_1r1w.synth.nz.mem[760] [12];
  assign _14101_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [12] : \MSYNC_1r1w.synth.nz.mem[762] [12];
  assign _14102_ = \bapg_rd.w_ptr_r [1] ? _14101_ : _14100_;
  assign _14103_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [12] : \MSYNC_1r1w.synth.nz.mem[764] [12];
  assign _14104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [12] : \MSYNC_1r1w.synth.nz.mem[766] [12];
  assign _14105_ = \bapg_rd.w_ptr_r [1] ? _14104_ : _14103_;
  assign _14106_ = \bapg_rd.w_ptr_r [2] ? _14105_ : _14102_;
  assign _14107_ = \bapg_rd.w_ptr_r [3] ? _14106_ : _14099_;
  assign _14108_ = \bapg_rd.w_ptr_r [4] ? _14107_ : _14092_;
  assign _14109_ = \bapg_rd.w_ptr_r [5] ? _14108_ : _14077_;
  assign _14110_ = \bapg_rd.w_ptr_r [6] ? _14109_ : _14046_;
  assign _14111_ = \bapg_rd.w_ptr_r [7] ? _14110_ : _13983_;
  assign _14112_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [12] : \MSYNC_1r1w.synth.nz.mem[768] [12];
  assign _14113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [12] : \MSYNC_1r1w.synth.nz.mem[770] [12];
  assign _14114_ = \bapg_rd.w_ptr_r [1] ? _14113_ : _14112_;
  assign _14115_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [12] : \MSYNC_1r1w.synth.nz.mem[772] [12];
  assign _14116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [12] : \MSYNC_1r1w.synth.nz.mem[774] [12];
  assign _14117_ = \bapg_rd.w_ptr_r [1] ? _14116_ : _14115_;
  assign _14118_ = \bapg_rd.w_ptr_r [2] ? _14117_ : _14114_;
  assign _14119_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [12] : \MSYNC_1r1w.synth.nz.mem[776] [12];
  assign _14120_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [12] : \MSYNC_1r1w.synth.nz.mem[778] [12];
  assign _14121_ = \bapg_rd.w_ptr_r [1] ? _14120_ : _14119_;
  assign _14122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [12] : \MSYNC_1r1w.synth.nz.mem[780] [12];
  assign _14123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [12] : \MSYNC_1r1w.synth.nz.mem[782] [12];
  assign _14124_ = \bapg_rd.w_ptr_r [1] ? _14123_ : _14122_;
  assign _14125_ = \bapg_rd.w_ptr_r [2] ? _14124_ : _14121_;
  assign _14126_ = \bapg_rd.w_ptr_r [3] ? _14125_ : _14118_;
  assign _14127_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [12] : \MSYNC_1r1w.synth.nz.mem[784] [12];
  assign _14128_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [12] : \MSYNC_1r1w.synth.nz.mem[786] [12];
  assign _14129_ = \bapg_rd.w_ptr_r [1] ? _14128_ : _14127_;
  assign _14130_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [12] : \MSYNC_1r1w.synth.nz.mem[788] [12];
  assign _14131_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [12] : \MSYNC_1r1w.synth.nz.mem[790] [12];
  assign _14132_ = \bapg_rd.w_ptr_r [1] ? _14131_ : _14130_;
  assign _14133_ = \bapg_rd.w_ptr_r [2] ? _14132_ : _14129_;
  assign _14134_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [12] : \MSYNC_1r1w.synth.nz.mem[792] [12];
  assign _14135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [12] : \MSYNC_1r1w.synth.nz.mem[794] [12];
  assign _14136_ = \bapg_rd.w_ptr_r [1] ? _14135_ : _14134_;
  assign _14137_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [12] : \MSYNC_1r1w.synth.nz.mem[796] [12];
  assign _14138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [12] : \MSYNC_1r1w.synth.nz.mem[798] [12];
  assign _14139_ = \bapg_rd.w_ptr_r [1] ? _14138_ : _14137_;
  assign _14140_ = \bapg_rd.w_ptr_r [2] ? _14139_ : _14136_;
  assign _14141_ = \bapg_rd.w_ptr_r [3] ? _14140_ : _14133_;
  assign _14142_ = \bapg_rd.w_ptr_r [4] ? _14141_ : _14126_;
  assign _14143_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [12] : \MSYNC_1r1w.synth.nz.mem[800] [12];
  assign _14144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [12] : \MSYNC_1r1w.synth.nz.mem[802] [12];
  assign _14145_ = \bapg_rd.w_ptr_r [1] ? _14144_ : _14143_;
  assign _14146_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [12] : \MSYNC_1r1w.synth.nz.mem[804] [12];
  assign _14147_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [12] : \MSYNC_1r1w.synth.nz.mem[806] [12];
  assign _14148_ = \bapg_rd.w_ptr_r [1] ? _14147_ : _14146_;
  assign _14149_ = \bapg_rd.w_ptr_r [2] ? _14148_ : _14145_;
  assign _14150_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [12] : \MSYNC_1r1w.synth.nz.mem[808] [12];
  assign _14151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [12] : \MSYNC_1r1w.synth.nz.mem[810] [12];
  assign _14152_ = \bapg_rd.w_ptr_r [1] ? _14151_ : _14150_;
  assign _14153_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [12] : \MSYNC_1r1w.synth.nz.mem[812] [12];
  assign _14154_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [12] : \MSYNC_1r1w.synth.nz.mem[814] [12];
  assign _14155_ = \bapg_rd.w_ptr_r [1] ? _14154_ : _14153_;
  assign _14156_ = \bapg_rd.w_ptr_r [2] ? _14155_ : _14152_;
  assign _14157_ = \bapg_rd.w_ptr_r [3] ? _14156_ : _14149_;
  assign _14158_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [12] : \MSYNC_1r1w.synth.nz.mem[816] [12];
  assign _14159_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [12] : \MSYNC_1r1w.synth.nz.mem[818] [12];
  assign _14160_ = \bapg_rd.w_ptr_r [1] ? _14159_ : _14158_;
  assign _14161_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [12] : \MSYNC_1r1w.synth.nz.mem[820] [12];
  assign _14162_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [12] : \MSYNC_1r1w.synth.nz.mem[822] [12];
  assign _14163_ = \bapg_rd.w_ptr_r [1] ? _14162_ : _14161_;
  assign _14164_ = \bapg_rd.w_ptr_r [2] ? _14163_ : _14160_;
  assign _14165_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [12] : \MSYNC_1r1w.synth.nz.mem[824] [12];
  assign _14166_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [12] : \MSYNC_1r1w.synth.nz.mem[826] [12];
  assign _14167_ = \bapg_rd.w_ptr_r [1] ? _14166_ : _14165_;
  assign _14168_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [12] : \MSYNC_1r1w.synth.nz.mem[828] [12];
  assign _14169_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [12] : \MSYNC_1r1w.synth.nz.mem[830] [12];
  assign _14170_ = \bapg_rd.w_ptr_r [1] ? _14169_ : _14168_;
  assign _14171_ = \bapg_rd.w_ptr_r [2] ? _14170_ : _14167_;
  assign _14172_ = \bapg_rd.w_ptr_r [3] ? _14171_ : _14164_;
  assign _14173_ = \bapg_rd.w_ptr_r [4] ? _14172_ : _14157_;
  assign _14174_ = \bapg_rd.w_ptr_r [5] ? _14173_ : _14142_;
  assign _14175_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [12] : \MSYNC_1r1w.synth.nz.mem[832] [12];
  assign _14176_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [12] : \MSYNC_1r1w.synth.nz.mem[834] [12];
  assign _14177_ = \bapg_rd.w_ptr_r [1] ? _14176_ : _14175_;
  assign _14178_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [12] : \MSYNC_1r1w.synth.nz.mem[836] [12];
  assign _14179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [12] : \MSYNC_1r1w.synth.nz.mem[838] [12];
  assign _14180_ = \bapg_rd.w_ptr_r [1] ? _14179_ : _14178_;
  assign _14181_ = \bapg_rd.w_ptr_r [2] ? _14180_ : _14177_;
  assign _14182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [12] : \MSYNC_1r1w.synth.nz.mem[840] [12];
  assign _14183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [12] : \MSYNC_1r1w.synth.nz.mem[842] [12];
  assign _14184_ = \bapg_rd.w_ptr_r [1] ? _14183_ : _14182_;
  assign _14185_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [12] : \MSYNC_1r1w.synth.nz.mem[844] [12];
  assign _14186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [12] : \MSYNC_1r1w.synth.nz.mem[846] [12];
  assign _14187_ = \bapg_rd.w_ptr_r [1] ? _14186_ : _14185_;
  assign _14188_ = \bapg_rd.w_ptr_r [2] ? _14187_ : _14184_;
  assign _14189_ = \bapg_rd.w_ptr_r [3] ? _14188_ : _14181_;
  assign _14190_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [12] : \MSYNC_1r1w.synth.nz.mem[848] [12];
  assign _14191_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [12] : \MSYNC_1r1w.synth.nz.mem[850] [12];
  assign _14192_ = \bapg_rd.w_ptr_r [1] ? _14191_ : _14190_;
  assign _14193_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [12] : \MSYNC_1r1w.synth.nz.mem[852] [12];
  assign _14194_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [12] : \MSYNC_1r1w.synth.nz.mem[854] [12];
  assign _14195_ = \bapg_rd.w_ptr_r [1] ? _14194_ : _14193_;
  assign _14196_ = \bapg_rd.w_ptr_r [2] ? _14195_ : _14192_;
  assign _14197_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [12] : \MSYNC_1r1w.synth.nz.mem[856] [12];
  assign _14198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [12] : \MSYNC_1r1w.synth.nz.mem[858] [12];
  assign _14199_ = \bapg_rd.w_ptr_r [1] ? _14198_ : _14197_;
  assign _14200_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [12] : \MSYNC_1r1w.synth.nz.mem[860] [12];
  assign _14201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [12] : \MSYNC_1r1w.synth.nz.mem[862] [12];
  assign _14202_ = \bapg_rd.w_ptr_r [1] ? _14201_ : _14200_;
  assign _14203_ = \bapg_rd.w_ptr_r [2] ? _14202_ : _14199_;
  assign _14204_ = \bapg_rd.w_ptr_r [3] ? _14203_ : _14196_;
  assign _14205_ = \bapg_rd.w_ptr_r [4] ? _14204_ : _14189_;
  assign _14206_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [12] : \MSYNC_1r1w.synth.nz.mem[864] [12];
  assign _14207_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [12] : \MSYNC_1r1w.synth.nz.mem[866] [12];
  assign _14208_ = \bapg_rd.w_ptr_r [1] ? _14207_ : _14206_;
  assign _14209_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [12] : \MSYNC_1r1w.synth.nz.mem[868] [12];
  assign _14210_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [12] : \MSYNC_1r1w.synth.nz.mem[870] [12];
  assign _14211_ = \bapg_rd.w_ptr_r [1] ? _14210_ : _14209_;
  assign _14212_ = \bapg_rd.w_ptr_r [2] ? _14211_ : _14208_;
  assign _14213_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [12] : \MSYNC_1r1w.synth.nz.mem[872] [12];
  assign _14214_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [12] : \MSYNC_1r1w.synth.nz.mem[874] [12];
  assign _14215_ = \bapg_rd.w_ptr_r [1] ? _14214_ : _14213_;
  assign _14216_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [12] : \MSYNC_1r1w.synth.nz.mem[876] [12];
  assign _14217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [12] : \MSYNC_1r1w.synth.nz.mem[878] [12];
  assign _14218_ = \bapg_rd.w_ptr_r [1] ? _14217_ : _14216_;
  assign _14219_ = \bapg_rd.w_ptr_r [2] ? _14218_ : _14215_;
  assign _14220_ = \bapg_rd.w_ptr_r [3] ? _14219_ : _14212_;
  assign _14221_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [12] : \MSYNC_1r1w.synth.nz.mem[880] [12];
  assign _14222_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [12] : \MSYNC_1r1w.synth.nz.mem[882] [12];
  assign _14223_ = \bapg_rd.w_ptr_r [1] ? _14222_ : _14221_;
  assign _14224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [12] : \MSYNC_1r1w.synth.nz.mem[884] [12];
  assign _14225_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [12] : \MSYNC_1r1w.synth.nz.mem[886] [12];
  assign _14226_ = \bapg_rd.w_ptr_r [1] ? _14225_ : _14224_;
  assign _14227_ = \bapg_rd.w_ptr_r [2] ? _14226_ : _14223_;
  assign _14228_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [12] : \MSYNC_1r1w.synth.nz.mem[888] [12];
  assign _14229_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [12] : \MSYNC_1r1w.synth.nz.mem[890] [12];
  assign _14230_ = \bapg_rd.w_ptr_r [1] ? _14229_ : _14228_;
  assign _14231_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [12] : \MSYNC_1r1w.synth.nz.mem[892] [12];
  assign _14232_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [12] : \MSYNC_1r1w.synth.nz.mem[894] [12];
  assign _14233_ = \bapg_rd.w_ptr_r [1] ? _14232_ : _14231_;
  assign _14234_ = \bapg_rd.w_ptr_r [2] ? _14233_ : _14230_;
  assign _14235_ = \bapg_rd.w_ptr_r [3] ? _14234_ : _14227_;
  assign _14236_ = \bapg_rd.w_ptr_r [4] ? _14235_ : _14220_;
  assign _14237_ = \bapg_rd.w_ptr_r [5] ? _14236_ : _14205_;
  assign _14238_ = \bapg_rd.w_ptr_r [6] ? _14237_ : _14174_;
  assign _14239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [12] : \MSYNC_1r1w.synth.nz.mem[896] [12];
  assign _14240_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [12] : \MSYNC_1r1w.synth.nz.mem[898] [12];
  assign _14241_ = \bapg_rd.w_ptr_r [1] ? _14240_ : _14239_;
  assign _14242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [12] : \MSYNC_1r1w.synth.nz.mem[900] [12];
  assign _14243_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [12] : \MSYNC_1r1w.synth.nz.mem[902] [12];
  assign _14244_ = \bapg_rd.w_ptr_r [1] ? _14243_ : _14242_;
  assign _14245_ = \bapg_rd.w_ptr_r [2] ? _14244_ : _14241_;
  assign _14246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [12] : \MSYNC_1r1w.synth.nz.mem[904] [12];
  assign _14247_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [12] : \MSYNC_1r1w.synth.nz.mem[906] [12];
  assign _14248_ = \bapg_rd.w_ptr_r [1] ? _14247_ : _14246_;
  assign _14249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [12] : \MSYNC_1r1w.synth.nz.mem[908] [12];
  assign _14250_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [12] : \MSYNC_1r1w.synth.nz.mem[910] [12];
  assign _14251_ = \bapg_rd.w_ptr_r [1] ? _14250_ : _14249_;
  assign _14252_ = \bapg_rd.w_ptr_r [2] ? _14251_ : _14248_;
  assign _14253_ = \bapg_rd.w_ptr_r [3] ? _14252_ : _14245_;
  assign _14254_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [12] : \MSYNC_1r1w.synth.nz.mem[912] [12];
  assign _14255_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [12] : \MSYNC_1r1w.synth.nz.mem[914] [12];
  assign _14256_ = \bapg_rd.w_ptr_r [1] ? _14255_ : _14254_;
  assign _14257_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [12] : \MSYNC_1r1w.synth.nz.mem[916] [12];
  assign _14258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [12] : \MSYNC_1r1w.synth.nz.mem[918] [12];
  assign _14259_ = \bapg_rd.w_ptr_r [1] ? _14258_ : _14257_;
  assign _14260_ = \bapg_rd.w_ptr_r [2] ? _14259_ : _14256_;
  assign _14261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [12] : \MSYNC_1r1w.synth.nz.mem[920] [12];
  assign _14262_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [12] : \MSYNC_1r1w.synth.nz.mem[922] [12];
  assign _14263_ = \bapg_rd.w_ptr_r [1] ? _14262_ : _14261_;
  assign _14264_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [12] : \MSYNC_1r1w.synth.nz.mem[924] [12];
  assign _14265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [12] : \MSYNC_1r1w.synth.nz.mem[926] [12];
  assign _14266_ = \bapg_rd.w_ptr_r [1] ? _14265_ : _14264_;
  assign _14267_ = \bapg_rd.w_ptr_r [2] ? _14266_ : _14263_;
  assign _14268_ = \bapg_rd.w_ptr_r [3] ? _14267_ : _14260_;
  assign _14269_ = \bapg_rd.w_ptr_r [4] ? _14268_ : _14253_;
  assign _14270_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [12] : \MSYNC_1r1w.synth.nz.mem[928] [12];
  assign _14271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [12] : \MSYNC_1r1w.synth.nz.mem[930] [12];
  assign _14272_ = \bapg_rd.w_ptr_r [1] ? _14271_ : _14270_;
  assign _14273_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [12] : \MSYNC_1r1w.synth.nz.mem[932] [12];
  assign _14274_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [12] : \MSYNC_1r1w.synth.nz.mem[934] [12];
  assign _14275_ = \bapg_rd.w_ptr_r [1] ? _14274_ : _14273_;
  assign _14276_ = \bapg_rd.w_ptr_r [2] ? _14275_ : _14272_;
  assign _14277_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [12] : \MSYNC_1r1w.synth.nz.mem[936] [12];
  assign _14278_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [12] : \MSYNC_1r1w.synth.nz.mem[938] [12];
  assign _14279_ = \bapg_rd.w_ptr_r [1] ? _14278_ : _14277_;
  assign _14280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [12] : \MSYNC_1r1w.synth.nz.mem[940] [12];
  assign _14281_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [12] : \MSYNC_1r1w.synth.nz.mem[942] [12];
  assign _14282_ = \bapg_rd.w_ptr_r [1] ? _14281_ : _14280_;
  assign _14283_ = \bapg_rd.w_ptr_r [2] ? _14282_ : _14279_;
  assign _14284_ = \bapg_rd.w_ptr_r [3] ? _14283_ : _14276_;
  assign _14285_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [12] : \MSYNC_1r1w.synth.nz.mem[944] [12];
  assign _14286_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [12] : \MSYNC_1r1w.synth.nz.mem[946] [12];
  assign _14287_ = \bapg_rd.w_ptr_r [1] ? _14286_ : _14285_;
  assign _14288_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [12] : \MSYNC_1r1w.synth.nz.mem[948] [12];
  assign _14289_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [12] : \MSYNC_1r1w.synth.nz.mem[950] [12];
  assign _14290_ = \bapg_rd.w_ptr_r [1] ? _14289_ : _14288_;
  assign _14291_ = \bapg_rd.w_ptr_r [2] ? _14290_ : _14287_;
  assign _14292_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [12] : \MSYNC_1r1w.synth.nz.mem[952] [12];
  assign _14293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [12] : \MSYNC_1r1w.synth.nz.mem[954] [12];
  assign _14294_ = \bapg_rd.w_ptr_r [1] ? _14293_ : _14292_;
  assign _14295_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [12] : \MSYNC_1r1w.synth.nz.mem[956] [12];
  assign _14296_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [12] : \MSYNC_1r1w.synth.nz.mem[958] [12];
  assign _14297_ = \bapg_rd.w_ptr_r [1] ? _14296_ : _14295_;
  assign _14298_ = \bapg_rd.w_ptr_r [2] ? _14297_ : _14294_;
  assign _14299_ = \bapg_rd.w_ptr_r [3] ? _14298_ : _14291_;
  assign _14300_ = \bapg_rd.w_ptr_r [4] ? _14299_ : _14284_;
  assign _14301_ = \bapg_rd.w_ptr_r [5] ? _14300_ : _14269_;
  assign _14302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [12] : \MSYNC_1r1w.synth.nz.mem[960] [12];
  assign _14303_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [12] : \MSYNC_1r1w.synth.nz.mem[962] [12];
  assign _14304_ = \bapg_rd.w_ptr_r [1] ? _14303_ : _14302_;
  assign _14305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [12] : \MSYNC_1r1w.synth.nz.mem[964] [12];
  assign _14306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [12] : \MSYNC_1r1w.synth.nz.mem[966] [12];
  assign _14307_ = \bapg_rd.w_ptr_r [1] ? _14306_ : _14305_;
  assign _14308_ = \bapg_rd.w_ptr_r [2] ? _14307_ : _14304_;
  assign _14309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [12] : \MSYNC_1r1w.synth.nz.mem[968] [12];
  assign _14310_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [12] : \MSYNC_1r1w.synth.nz.mem[970] [12];
  assign _14311_ = \bapg_rd.w_ptr_r [1] ? _14310_ : _14309_;
  assign _14312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [12] : \MSYNC_1r1w.synth.nz.mem[972] [12];
  assign _14313_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [12] : \MSYNC_1r1w.synth.nz.mem[974] [12];
  assign _14314_ = \bapg_rd.w_ptr_r [1] ? _14313_ : _14312_;
  assign _14315_ = \bapg_rd.w_ptr_r [2] ? _14314_ : _14311_;
  assign _14316_ = \bapg_rd.w_ptr_r [3] ? _14315_ : _14308_;
  assign _14317_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [12] : \MSYNC_1r1w.synth.nz.mem[976] [12];
  assign _14318_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [12] : \MSYNC_1r1w.synth.nz.mem[978] [12];
  assign _14319_ = \bapg_rd.w_ptr_r [1] ? _14318_ : _14317_;
  assign _14320_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [12] : \MSYNC_1r1w.synth.nz.mem[980] [12];
  assign _14321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [12] : \MSYNC_1r1w.synth.nz.mem[982] [12];
  assign _14322_ = \bapg_rd.w_ptr_r [1] ? _14321_ : _14320_;
  assign _14323_ = \bapg_rd.w_ptr_r [2] ? _14322_ : _14319_;
  assign _14324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [12] : \MSYNC_1r1w.synth.nz.mem[984] [12];
  assign _14325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [12] : \MSYNC_1r1w.synth.nz.mem[986] [12];
  assign _14326_ = \bapg_rd.w_ptr_r [1] ? _14325_ : _14324_;
  assign _14327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [12] : \MSYNC_1r1w.synth.nz.mem[988] [12];
  assign _14328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [12] : \MSYNC_1r1w.synth.nz.mem[990] [12];
  assign _14329_ = \bapg_rd.w_ptr_r [1] ? _14328_ : _14327_;
  assign _14330_ = \bapg_rd.w_ptr_r [2] ? _14329_ : _14326_;
  assign _14331_ = \bapg_rd.w_ptr_r [3] ? _14330_ : _14323_;
  assign _14332_ = \bapg_rd.w_ptr_r [4] ? _14331_ : _14316_;
  assign _14333_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [12] : \MSYNC_1r1w.synth.nz.mem[992] [12];
  assign _14334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [12] : \MSYNC_1r1w.synth.nz.mem[994] [12];
  assign _14335_ = \bapg_rd.w_ptr_r [1] ? _14334_ : _14333_;
  assign _14336_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [12] : \MSYNC_1r1w.synth.nz.mem[996] [12];
  assign _14337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [12] : \MSYNC_1r1w.synth.nz.mem[998] [12];
  assign _14338_ = \bapg_rd.w_ptr_r [1] ? _14337_ : _14336_;
  assign _14339_ = \bapg_rd.w_ptr_r [2] ? _14338_ : _14335_;
  assign _14340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [12] : \MSYNC_1r1w.synth.nz.mem[1000] [12];
  assign _14341_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [12] : \MSYNC_1r1w.synth.nz.mem[1002] [12];
  assign _14342_ = \bapg_rd.w_ptr_r [1] ? _14341_ : _14340_;
  assign _14343_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [12] : \MSYNC_1r1w.synth.nz.mem[1004] [12];
  assign _14344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [12] : \MSYNC_1r1w.synth.nz.mem[1006] [12];
  assign _14345_ = \bapg_rd.w_ptr_r [1] ? _14344_ : _14343_;
  assign _14346_ = \bapg_rd.w_ptr_r [2] ? _14345_ : _14342_;
  assign _14347_ = \bapg_rd.w_ptr_r [3] ? _14346_ : _14339_;
  assign _14348_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [12] : \MSYNC_1r1w.synth.nz.mem[1008] [12];
  assign _14349_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [12] : \MSYNC_1r1w.synth.nz.mem[1010] [12];
  assign _14350_ = \bapg_rd.w_ptr_r [1] ? _14349_ : _14348_;
  assign _14351_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [12] : \MSYNC_1r1w.synth.nz.mem[1012] [12];
  assign _14352_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [12] : \MSYNC_1r1w.synth.nz.mem[1014] [12];
  assign _14353_ = \bapg_rd.w_ptr_r [1] ? _14352_ : _14351_;
  assign _14354_ = \bapg_rd.w_ptr_r [2] ? _14353_ : _14350_;
  assign _14355_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [12] : \MSYNC_1r1w.synth.nz.mem[1016] [12];
  assign _14356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [12] : \MSYNC_1r1w.synth.nz.mem[1018] [12];
  assign _14357_ = \bapg_rd.w_ptr_r [1] ? _14356_ : _14355_;
  assign _14358_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [12] : \MSYNC_1r1w.synth.nz.mem[1020] [12];
  assign _14359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [12] : \MSYNC_1r1w.synth.nz.mem[1022] [12];
  assign _14360_ = \bapg_rd.w_ptr_r [1] ? _14359_ : _14358_;
  assign _14361_ = \bapg_rd.w_ptr_r [2] ? _14360_ : _14357_;
  assign _14362_ = \bapg_rd.w_ptr_r [3] ? _14361_ : _14354_;
  assign _14363_ = \bapg_rd.w_ptr_r [4] ? _14362_ : _14347_;
  assign _14364_ = \bapg_rd.w_ptr_r [5] ? _14363_ : _14332_;
  assign _14365_ = \bapg_rd.w_ptr_r [6] ? _14364_ : _14301_;
  assign _14366_ = \bapg_rd.w_ptr_r [7] ? _14365_ : _14238_;
  assign _14367_ = \bapg_rd.w_ptr_r [8] ? _14366_ : _14111_;
  assign r_data_o[12] = \bapg_rd.w_ptr_r [9] ? _14367_ : _13856_;
  assign _14368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [13] : \MSYNC_1r1w.synth.nz.mem[0] [13];
  assign _14369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [13] : \MSYNC_1r1w.synth.nz.mem[2] [13];
  assign _14370_ = \bapg_rd.w_ptr_r [1] ? _14369_ : _14368_;
  assign _14371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [13] : \MSYNC_1r1w.synth.nz.mem[4] [13];
  assign _14372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [13] : \MSYNC_1r1w.synth.nz.mem[6] [13];
  assign _14373_ = \bapg_rd.w_ptr_r [1] ? _14372_ : _14371_;
  assign _14374_ = \bapg_rd.w_ptr_r [2] ? _14373_ : _14370_;
  assign _14375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [13] : \MSYNC_1r1w.synth.nz.mem[8] [13];
  assign _14376_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [13] : \MSYNC_1r1w.synth.nz.mem[10] [13];
  assign _14377_ = \bapg_rd.w_ptr_r [1] ? _14376_ : _14375_;
  assign _14378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [13] : \MSYNC_1r1w.synth.nz.mem[12] [13];
  assign _14379_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [13] : \MSYNC_1r1w.synth.nz.mem[14] [13];
  assign _14380_ = \bapg_rd.w_ptr_r [1] ? _14379_ : _14378_;
  assign _14381_ = \bapg_rd.w_ptr_r [2] ? _14380_ : _14377_;
  assign _14382_ = \bapg_rd.w_ptr_r [3] ? _14381_ : _14374_;
  assign _14383_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [13] : \MSYNC_1r1w.synth.nz.mem[16] [13];
  assign _14384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [13] : \MSYNC_1r1w.synth.nz.mem[18] [13];
  assign _14385_ = \bapg_rd.w_ptr_r [1] ? _14384_ : _14383_;
  assign _14386_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [13] : \MSYNC_1r1w.synth.nz.mem[20] [13];
  assign _14387_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [13] : \MSYNC_1r1w.synth.nz.mem[22] [13];
  assign _14388_ = \bapg_rd.w_ptr_r [1] ? _14387_ : _14386_;
  assign _14389_ = \bapg_rd.w_ptr_r [2] ? _14388_ : _14385_;
  assign _14390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [13] : \MSYNC_1r1w.synth.nz.mem[24] [13];
  assign _14391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [13] : \MSYNC_1r1w.synth.nz.mem[26] [13];
  assign _14392_ = \bapg_rd.w_ptr_r [1] ? _14391_ : _14390_;
  assign _14393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [13] : \MSYNC_1r1w.synth.nz.mem[28] [13];
  assign _14394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [13] : \MSYNC_1r1w.synth.nz.mem[30] [13];
  assign _14395_ = \bapg_rd.w_ptr_r [1] ? _14394_ : _14393_;
  assign _14396_ = \bapg_rd.w_ptr_r [2] ? _14395_ : _14392_;
  assign _14397_ = \bapg_rd.w_ptr_r [3] ? _14396_ : _14389_;
  assign _14398_ = \bapg_rd.w_ptr_r [4] ? _14397_ : _14382_;
  assign _14399_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [13] : \MSYNC_1r1w.synth.nz.mem[32] [13];
  assign _14400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [13] : \MSYNC_1r1w.synth.nz.mem[34] [13];
  assign _14401_ = \bapg_rd.w_ptr_r [1] ? _14400_ : _14399_;
  assign _14402_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [13] : \MSYNC_1r1w.synth.nz.mem[36] [13];
  assign _14403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [13] : \MSYNC_1r1w.synth.nz.mem[38] [13];
  assign _14404_ = \bapg_rd.w_ptr_r [1] ? _14403_ : _14402_;
  assign _14405_ = \bapg_rd.w_ptr_r [2] ? _14404_ : _14401_;
  assign _14406_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [13] : \MSYNC_1r1w.synth.nz.mem[40] [13];
  assign _14407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [13] : \MSYNC_1r1w.synth.nz.mem[42] [13];
  assign _14408_ = \bapg_rd.w_ptr_r [1] ? _14407_ : _14406_;
  assign _14409_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [13] : \MSYNC_1r1w.synth.nz.mem[44] [13];
  assign _14410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [13] : \MSYNC_1r1w.synth.nz.mem[46] [13];
  assign _14411_ = \bapg_rd.w_ptr_r [1] ? _14410_ : _14409_;
  assign _14412_ = \bapg_rd.w_ptr_r [2] ? _14411_ : _14408_;
  assign _14413_ = \bapg_rd.w_ptr_r [3] ? _14412_ : _14405_;
  assign _14414_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [13] : \MSYNC_1r1w.synth.nz.mem[48] [13];
  assign _14415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [13] : \MSYNC_1r1w.synth.nz.mem[50] [13];
  assign _14416_ = \bapg_rd.w_ptr_r [1] ? _14415_ : _14414_;
  assign _14417_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [13] : \MSYNC_1r1w.synth.nz.mem[52] [13];
  assign _14418_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [13] : \MSYNC_1r1w.synth.nz.mem[54] [13];
  assign _14419_ = \bapg_rd.w_ptr_r [1] ? _14418_ : _14417_;
  assign _14420_ = \bapg_rd.w_ptr_r [2] ? _14419_ : _14416_;
  assign _14421_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [13] : \MSYNC_1r1w.synth.nz.mem[56] [13];
  assign _14422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [13] : \MSYNC_1r1w.synth.nz.mem[58] [13];
  assign _14423_ = \bapg_rd.w_ptr_r [1] ? _14422_ : _14421_;
  assign _14424_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [13] : \MSYNC_1r1w.synth.nz.mem[60] [13];
  assign _14425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [13] : \MSYNC_1r1w.synth.nz.mem[62] [13];
  assign _14426_ = \bapg_rd.w_ptr_r [1] ? _14425_ : _14424_;
  assign _14427_ = \bapg_rd.w_ptr_r [2] ? _14426_ : _14423_;
  assign _14428_ = \bapg_rd.w_ptr_r [3] ? _14427_ : _14420_;
  assign _14429_ = \bapg_rd.w_ptr_r [4] ? _14428_ : _14413_;
  assign _14430_ = \bapg_rd.w_ptr_r [5] ? _14429_ : _14398_;
  assign _14431_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [13] : \MSYNC_1r1w.synth.nz.mem[64] [13];
  assign _14432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [13] : \MSYNC_1r1w.synth.nz.mem[66] [13];
  assign _14433_ = \bapg_rd.w_ptr_r [1] ? _14432_ : _14431_;
  assign _14434_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [13] : \MSYNC_1r1w.synth.nz.mem[68] [13];
  assign _14435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [13] : \MSYNC_1r1w.synth.nz.mem[70] [13];
  assign _14436_ = \bapg_rd.w_ptr_r [1] ? _14435_ : _14434_;
  assign _14437_ = \bapg_rd.w_ptr_r [2] ? _14436_ : _14433_;
  assign _14438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [13] : \MSYNC_1r1w.synth.nz.mem[72] [13];
  assign _14439_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [13] : \MSYNC_1r1w.synth.nz.mem[74] [13];
  assign _14440_ = \bapg_rd.w_ptr_r [1] ? _14439_ : _14438_;
  assign _14441_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [13] : \MSYNC_1r1w.synth.nz.mem[76] [13];
  assign _14442_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [13] : \MSYNC_1r1w.synth.nz.mem[78] [13];
  assign _14443_ = \bapg_rd.w_ptr_r [1] ? _14442_ : _14441_;
  assign _14444_ = \bapg_rd.w_ptr_r [2] ? _14443_ : _14440_;
  assign _14445_ = \bapg_rd.w_ptr_r [3] ? _14444_ : _14437_;
  assign _14446_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [13] : \MSYNC_1r1w.synth.nz.mem[80] [13];
  assign _14447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [13] : \MSYNC_1r1w.synth.nz.mem[82] [13];
  assign _14448_ = \bapg_rd.w_ptr_r [1] ? _14447_ : _14446_;
  assign _14449_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [13] : \MSYNC_1r1w.synth.nz.mem[84] [13];
  assign _14450_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [13] : \MSYNC_1r1w.synth.nz.mem[86] [13];
  assign _14451_ = \bapg_rd.w_ptr_r [1] ? _14450_ : _14449_;
  assign _14452_ = \bapg_rd.w_ptr_r [2] ? _14451_ : _14448_;
  assign _14453_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [13] : \MSYNC_1r1w.synth.nz.mem[88] [13];
  assign _14454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [13] : \MSYNC_1r1w.synth.nz.mem[90] [13];
  assign _14455_ = \bapg_rd.w_ptr_r [1] ? _14454_ : _14453_;
  assign _14456_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [13] : \MSYNC_1r1w.synth.nz.mem[92] [13];
  assign _14457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [13] : \MSYNC_1r1w.synth.nz.mem[94] [13];
  assign _14458_ = \bapg_rd.w_ptr_r [1] ? _14457_ : _14456_;
  assign _14459_ = \bapg_rd.w_ptr_r [2] ? _14458_ : _14455_;
  assign _14460_ = \bapg_rd.w_ptr_r [3] ? _14459_ : _14452_;
  assign _14461_ = \bapg_rd.w_ptr_r [4] ? _14460_ : _14445_;
  assign _14462_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [13] : \MSYNC_1r1w.synth.nz.mem[96] [13];
  assign _14463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [13] : \MSYNC_1r1w.synth.nz.mem[98] [13];
  assign _14464_ = \bapg_rd.w_ptr_r [1] ? _14463_ : _14462_;
  assign _14465_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [13] : \MSYNC_1r1w.synth.nz.mem[100] [13];
  assign _14466_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [13] : \MSYNC_1r1w.synth.nz.mem[102] [13];
  assign _14467_ = \bapg_rd.w_ptr_r [1] ? _14466_ : _14465_;
  assign _14468_ = \bapg_rd.w_ptr_r [2] ? _14467_ : _14464_;
  assign _14469_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [13] : \MSYNC_1r1w.synth.nz.mem[104] [13];
  assign _14470_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [13] : \MSYNC_1r1w.synth.nz.mem[106] [13];
  assign _14471_ = \bapg_rd.w_ptr_r [1] ? _14470_ : _14469_;
  assign _14472_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [13] : \MSYNC_1r1w.synth.nz.mem[108] [13];
  assign _14473_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [13] : \MSYNC_1r1w.synth.nz.mem[110] [13];
  assign _14474_ = \bapg_rd.w_ptr_r [1] ? _14473_ : _14472_;
  assign _14475_ = \bapg_rd.w_ptr_r [2] ? _14474_ : _14471_;
  assign _14476_ = \bapg_rd.w_ptr_r [3] ? _14475_ : _14468_;
  assign _14477_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [13] : \MSYNC_1r1w.synth.nz.mem[112] [13];
  assign _14478_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [13] : \MSYNC_1r1w.synth.nz.mem[114] [13];
  assign _14479_ = \bapg_rd.w_ptr_r [1] ? _14478_ : _14477_;
  assign _14480_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [13] : \MSYNC_1r1w.synth.nz.mem[116] [13];
  assign _14481_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [13] : \MSYNC_1r1w.synth.nz.mem[118] [13];
  assign _14482_ = \bapg_rd.w_ptr_r [1] ? _14481_ : _14480_;
  assign _14483_ = \bapg_rd.w_ptr_r [2] ? _14482_ : _14479_;
  assign _14484_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [13] : \MSYNC_1r1w.synth.nz.mem[120] [13];
  assign _14485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [13] : \MSYNC_1r1w.synth.nz.mem[122] [13];
  assign _14486_ = \bapg_rd.w_ptr_r [1] ? _14485_ : _14484_;
  assign _14487_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [13] : \MSYNC_1r1w.synth.nz.mem[124] [13];
  assign _14488_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [13] : \MSYNC_1r1w.synth.nz.mem[126] [13];
  assign _14489_ = \bapg_rd.w_ptr_r [1] ? _14488_ : _14487_;
  assign _14490_ = \bapg_rd.w_ptr_r [2] ? _14489_ : _14486_;
  assign _14491_ = \bapg_rd.w_ptr_r [3] ? _14490_ : _14483_;
  assign _14492_ = \bapg_rd.w_ptr_r [4] ? _14491_ : _14476_;
  assign _14493_ = \bapg_rd.w_ptr_r [5] ? _14492_ : _14461_;
  assign _14494_ = \bapg_rd.w_ptr_r [6] ? _14493_ : _14430_;
  assign _14495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [13] : \MSYNC_1r1w.synth.nz.mem[128] [13];
  assign _14496_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [13] : \MSYNC_1r1w.synth.nz.mem[130] [13];
  assign _14497_ = \bapg_rd.w_ptr_r [1] ? _14496_ : _14495_;
  assign _14498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [13] : \MSYNC_1r1w.synth.nz.mem[132] [13];
  assign _14499_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [13] : \MSYNC_1r1w.synth.nz.mem[134] [13];
  assign _14500_ = \bapg_rd.w_ptr_r [1] ? _14499_ : _14498_;
  assign _14501_ = \bapg_rd.w_ptr_r [2] ? _14500_ : _14497_;
  assign _14502_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [13] : \MSYNC_1r1w.synth.nz.mem[136] [13];
  assign _14503_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [13] : \MSYNC_1r1w.synth.nz.mem[138] [13];
  assign _14504_ = \bapg_rd.w_ptr_r [1] ? _14503_ : _14502_;
  assign _14505_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [13] : \MSYNC_1r1w.synth.nz.mem[140] [13];
  assign _14506_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [13] : \MSYNC_1r1w.synth.nz.mem[142] [13];
  assign _14507_ = \bapg_rd.w_ptr_r [1] ? _14506_ : _14505_;
  assign _14508_ = \bapg_rd.w_ptr_r [2] ? _14507_ : _14504_;
  assign _14509_ = \bapg_rd.w_ptr_r [3] ? _14508_ : _14501_;
  assign _14510_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [13] : \MSYNC_1r1w.synth.nz.mem[144] [13];
  assign _14511_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [13] : \MSYNC_1r1w.synth.nz.mem[146] [13];
  assign _14512_ = \bapg_rd.w_ptr_r [1] ? _14511_ : _14510_;
  assign _14513_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [13] : \MSYNC_1r1w.synth.nz.mem[148] [13];
  assign _14514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [13] : \MSYNC_1r1w.synth.nz.mem[150] [13];
  assign _14515_ = \bapg_rd.w_ptr_r [1] ? _14514_ : _14513_;
  assign _14516_ = \bapg_rd.w_ptr_r [2] ? _14515_ : _14512_;
  assign _14517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [13] : \MSYNC_1r1w.synth.nz.mem[152] [13];
  assign _14518_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [13] : \MSYNC_1r1w.synth.nz.mem[154] [13];
  assign _14519_ = \bapg_rd.w_ptr_r [1] ? _14518_ : _14517_;
  assign _14520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [13] : \MSYNC_1r1w.synth.nz.mem[156] [13];
  assign _14521_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [13] : \MSYNC_1r1w.synth.nz.mem[158] [13];
  assign _14522_ = \bapg_rd.w_ptr_r [1] ? _14521_ : _14520_;
  assign _14523_ = \bapg_rd.w_ptr_r [2] ? _14522_ : _14519_;
  assign _14524_ = \bapg_rd.w_ptr_r [3] ? _14523_ : _14516_;
  assign _14525_ = \bapg_rd.w_ptr_r [4] ? _14524_ : _14509_;
  assign _14526_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [13] : \MSYNC_1r1w.synth.nz.mem[160] [13];
  assign _14527_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [13] : \MSYNC_1r1w.synth.nz.mem[162] [13];
  assign _14528_ = \bapg_rd.w_ptr_r [1] ? _14527_ : _14526_;
  assign _14529_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [13] : \MSYNC_1r1w.synth.nz.mem[164] [13];
  assign _14530_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [13] : \MSYNC_1r1w.synth.nz.mem[166] [13];
  assign _14531_ = \bapg_rd.w_ptr_r [1] ? _14530_ : _14529_;
  assign _14532_ = \bapg_rd.w_ptr_r [2] ? _14531_ : _14528_;
  assign _14533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [13] : \MSYNC_1r1w.synth.nz.mem[168] [13];
  assign _14534_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [13] : \MSYNC_1r1w.synth.nz.mem[170] [13];
  assign _14535_ = \bapg_rd.w_ptr_r [1] ? _14534_ : _14533_;
  assign _14536_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [13] : \MSYNC_1r1w.synth.nz.mem[172] [13];
  assign _14537_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [13] : \MSYNC_1r1w.synth.nz.mem[174] [13];
  assign _14538_ = \bapg_rd.w_ptr_r [1] ? _14537_ : _14536_;
  assign _14539_ = \bapg_rd.w_ptr_r [2] ? _14538_ : _14535_;
  assign _14540_ = \bapg_rd.w_ptr_r [3] ? _14539_ : _14532_;
  assign _14541_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [13] : \MSYNC_1r1w.synth.nz.mem[176] [13];
  assign _14542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [13] : \MSYNC_1r1w.synth.nz.mem[178] [13];
  assign _14543_ = \bapg_rd.w_ptr_r [1] ? _14542_ : _14541_;
  assign _14544_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [13] : \MSYNC_1r1w.synth.nz.mem[180] [13];
  assign _14545_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [13] : \MSYNC_1r1w.synth.nz.mem[182] [13];
  assign _14546_ = \bapg_rd.w_ptr_r [1] ? _14545_ : _14544_;
  assign _14547_ = \bapg_rd.w_ptr_r [2] ? _14546_ : _14543_;
  assign _14548_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [13] : \MSYNC_1r1w.synth.nz.mem[184] [13];
  assign _14549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [13] : \MSYNC_1r1w.synth.nz.mem[186] [13];
  assign _14550_ = \bapg_rd.w_ptr_r [1] ? _14549_ : _14548_;
  assign _14551_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [13] : \MSYNC_1r1w.synth.nz.mem[188] [13];
  assign _14552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [13] : \MSYNC_1r1w.synth.nz.mem[190] [13];
  assign _14553_ = \bapg_rd.w_ptr_r [1] ? _14552_ : _14551_;
  assign _14554_ = \bapg_rd.w_ptr_r [2] ? _14553_ : _14550_;
  assign _14555_ = \bapg_rd.w_ptr_r [3] ? _14554_ : _14547_;
  assign _14556_ = \bapg_rd.w_ptr_r [4] ? _14555_ : _14540_;
  assign _14557_ = \bapg_rd.w_ptr_r [5] ? _14556_ : _14525_;
  assign _14558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [13] : \MSYNC_1r1w.synth.nz.mem[192] [13];
  assign _14559_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [13] : \MSYNC_1r1w.synth.nz.mem[194] [13];
  assign _14560_ = \bapg_rd.w_ptr_r [1] ? _14559_ : _14558_;
  assign _14561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [13] : \MSYNC_1r1w.synth.nz.mem[196] [13];
  assign _14562_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [13] : \MSYNC_1r1w.synth.nz.mem[198] [13];
  assign _14563_ = \bapg_rd.w_ptr_r [1] ? _14562_ : _14561_;
  assign _14564_ = \bapg_rd.w_ptr_r [2] ? _14563_ : _14560_;
  assign _14565_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [13] : \MSYNC_1r1w.synth.nz.mem[200] [13];
  assign _14566_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [13] : \MSYNC_1r1w.synth.nz.mem[202] [13];
  assign _14567_ = \bapg_rd.w_ptr_r [1] ? _14566_ : _14565_;
  assign _14568_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [13] : \MSYNC_1r1w.synth.nz.mem[204] [13];
  assign _14569_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [13] : \MSYNC_1r1w.synth.nz.mem[206] [13];
  assign _14570_ = \bapg_rd.w_ptr_r [1] ? _14569_ : _14568_;
  assign _14571_ = \bapg_rd.w_ptr_r [2] ? _14570_ : _14567_;
  assign _14572_ = \bapg_rd.w_ptr_r [3] ? _14571_ : _14564_;
  assign _14573_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [13] : \MSYNC_1r1w.synth.nz.mem[208] [13];
  assign _14574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [13] : \MSYNC_1r1w.synth.nz.mem[210] [13];
  assign _14575_ = \bapg_rd.w_ptr_r [1] ? _14574_ : _14573_;
  assign _14576_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [13] : \MSYNC_1r1w.synth.nz.mem[212] [13];
  assign _14577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [13] : \MSYNC_1r1w.synth.nz.mem[214] [13];
  assign _14578_ = \bapg_rd.w_ptr_r [1] ? _14577_ : _14576_;
  assign _14579_ = \bapg_rd.w_ptr_r [2] ? _14578_ : _14575_;
  assign _14580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [13] : \MSYNC_1r1w.synth.nz.mem[216] [13];
  assign _14581_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [13] : \MSYNC_1r1w.synth.nz.mem[218] [13];
  assign _14582_ = \bapg_rd.w_ptr_r [1] ? _14581_ : _14580_;
  assign _14583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [13] : \MSYNC_1r1w.synth.nz.mem[220] [13];
  assign _14584_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [13] : \MSYNC_1r1w.synth.nz.mem[222] [13];
  assign _14585_ = \bapg_rd.w_ptr_r [1] ? _14584_ : _14583_;
  assign _14586_ = \bapg_rd.w_ptr_r [2] ? _14585_ : _14582_;
  assign _14587_ = \bapg_rd.w_ptr_r [3] ? _14586_ : _14579_;
  assign _14588_ = \bapg_rd.w_ptr_r [4] ? _14587_ : _14572_;
  assign _14589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [13] : \MSYNC_1r1w.synth.nz.mem[224] [13];
  assign _14590_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [13] : \MSYNC_1r1w.synth.nz.mem[226] [13];
  assign _14591_ = \bapg_rd.w_ptr_r [1] ? _14590_ : _14589_;
  assign _14592_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [13] : \MSYNC_1r1w.synth.nz.mem[228] [13];
  assign _14593_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [13] : \MSYNC_1r1w.synth.nz.mem[230] [13];
  assign _14594_ = \bapg_rd.w_ptr_r [1] ? _14593_ : _14592_;
  assign _14595_ = \bapg_rd.w_ptr_r [2] ? _14594_ : _14591_;
  assign _14596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [13] : \MSYNC_1r1w.synth.nz.mem[232] [13];
  assign _14597_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [13] : \MSYNC_1r1w.synth.nz.mem[234] [13];
  assign _14598_ = \bapg_rd.w_ptr_r [1] ? _14597_ : _14596_;
  assign _14599_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [13] : \MSYNC_1r1w.synth.nz.mem[236] [13];
  assign _14600_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [13] : \MSYNC_1r1w.synth.nz.mem[238] [13];
  assign _14601_ = \bapg_rd.w_ptr_r [1] ? _14600_ : _14599_;
  assign _14602_ = \bapg_rd.w_ptr_r [2] ? _14601_ : _14598_;
  assign _14603_ = \bapg_rd.w_ptr_r [3] ? _14602_ : _14595_;
  assign _14604_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [13] : \MSYNC_1r1w.synth.nz.mem[240] [13];
  assign _14605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [13] : \MSYNC_1r1w.synth.nz.mem[242] [13];
  assign _14606_ = \bapg_rd.w_ptr_r [1] ? _14605_ : _14604_;
  assign _14607_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [13] : \MSYNC_1r1w.synth.nz.mem[244] [13];
  assign _14608_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [13] : \MSYNC_1r1w.synth.nz.mem[246] [13];
  assign _14609_ = \bapg_rd.w_ptr_r [1] ? _14608_ : _14607_;
  assign _14610_ = \bapg_rd.w_ptr_r [2] ? _14609_ : _14606_;
  assign _14611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [13] : \MSYNC_1r1w.synth.nz.mem[248] [13];
  assign _14612_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [13] : \MSYNC_1r1w.synth.nz.mem[250] [13];
  assign _14613_ = \bapg_rd.w_ptr_r [1] ? _14612_ : _14611_;
  assign _14614_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [13] : \MSYNC_1r1w.synth.nz.mem[252] [13];
  assign _14615_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [13] : \MSYNC_1r1w.synth.nz.mem[254] [13];
  assign _14616_ = \bapg_rd.w_ptr_r [1] ? _14615_ : _14614_;
  assign _14617_ = \bapg_rd.w_ptr_r [2] ? _14616_ : _14613_;
  assign _14618_ = \bapg_rd.w_ptr_r [3] ? _14617_ : _14610_;
  assign _14619_ = \bapg_rd.w_ptr_r [4] ? _14618_ : _14603_;
  assign _14620_ = \bapg_rd.w_ptr_r [5] ? _14619_ : _14588_;
  assign _14621_ = \bapg_rd.w_ptr_r [6] ? _14620_ : _14557_;
  assign _14622_ = \bapg_rd.w_ptr_r [7] ? _14621_ : _14494_;
  assign _14623_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [13] : \MSYNC_1r1w.synth.nz.mem[256] [13];
  assign _14624_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [13] : \MSYNC_1r1w.synth.nz.mem[258] [13];
  assign _14625_ = \bapg_rd.w_ptr_r [1] ? _14624_ : _14623_;
  assign _14626_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [13] : \MSYNC_1r1w.synth.nz.mem[260] [13];
  assign _14627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [13] : \MSYNC_1r1w.synth.nz.mem[262] [13];
  assign _14628_ = \bapg_rd.w_ptr_r [1] ? _14627_ : _14626_;
  assign _14629_ = \bapg_rd.w_ptr_r [2] ? _14628_ : _14625_;
  assign _14630_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [13] : \MSYNC_1r1w.synth.nz.mem[264] [13];
  assign _14631_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [13] : \MSYNC_1r1w.synth.nz.mem[266] [13];
  assign _14632_ = \bapg_rd.w_ptr_r [1] ? _14631_ : _14630_;
  assign _14633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [13] : \MSYNC_1r1w.synth.nz.mem[268] [13];
  assign _14634_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [13] : \MSYNC_1r1w.synth.nz.mem[270] [13];
  assign _14635_ = \bapg_rd.w_ptr_r [1] ? _14634_ : _14633_;
  assign _14636_ = \bapg_rd.w_ptr_r [2] ? _14635_ : _14632_;
  assign _14637_ = \bapg_rd.w_ptr_r [3] ? _14636_ : _14629_;
  assign _14638_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [13] : \MSYNC_1r1w.synth.nz.mem[272] [13];
  assign _14639_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [13] : \MSYNC_1r1w.synth.nz.mem[274] [13];
  assign _14640_ = \bapg_rd.w_ptr_r [1] ? _14639_ : _14638_;
  assign _14641_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [13] : \MSYNC_1r1w.synth.nz.mem[276] [13];
  assign _14642_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [13] : \MSYNC_1r1w.synth.nz.mem[278] [13];
  assign _14643_ = \bapg_rd.w_ptr_r [1] ? _14642_ : _14641_;
  assign _14644_ = \bapg_rd.w_ptr_r [2] ? _14643_ : _14640_;
  assign _14645_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [13] : \MSYNC_1r1w.synth.nz.mem[280] [13];
  assign _14646_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [13] : \MSYNC_1r1w.synth.nz.mem[282] [13];
  assign _14647_ = \bapg_rd.w_ptr_r [1] ? _14646_ : _14645_;
  assign _14648_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [13] : \MSYNC_1r1w.synth.nz.mem[284] [13];
  assign _14649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [13] : \MSYNC_1r1w.synth.nz.mem[286] [13];
  assign _14650_ = \bapg_rd.w_ptr_r [1] ? _14649_ : _14648_;
  assign _14651_ = \bapg_rd.w_ptr_r [2] ? _14650_ : _14647_;
  assign _14652_ = \bapg_rd.w_ptr_r [3] ? _14651_ : _14644_;
  assign _14653_ = \bapg_rd.w_ptr_r [4] ? _14652_ : _14637_;
  assign _14654_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [13] : \MSYNC_1r1w.synth.nz.mem[288] [13];
  assign _14655_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [13] : \MSYNC_1r1w.synth.nz.mem[290] [13];
  assign _14656_ = \bapg_rd.w_ptr_r [1] ? _14655_ : _14654_;
  assign _14657_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [13] : \MSYNC_1r1w.synth.nz.mem[292] [13];
  assign _14658_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [13] : \MSYNC_1r1w.synth.nz.mem[294] [13];
  assign _14659_ = \bapg_rd.w_ptr_r [1] ? _14658_ : _14657_;
  assign _14660_ = \bapg_rd.w_ptr_r [2] ? _14659_ : _14656_;
  assign _14661_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [13] : \MSYNC_1r1w.synth.nz.mem[296] [13];
  assign _14662_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [13] : \MSYNC_1r1w.synth.nz.mem[298] [13];
  assign _14663_ = \bapg_rd.w_ptr_r [1] ? _14662_ : _14661_;
  assign _14664_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [13] : \MSYNC_1r1w.synth.nz.mem[300] [13];
  assign _14665_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [13] : \MSYNC_1r1w.synth.nz.mem[302] [13];
  assign _14666_ = \bapg_rd.w_ptr_r [1] ? _14665_ : _14664_;
  assign _14667_ = \bapg_rd.w_ptr_r [2] ? _14666_ : _14663_;
  assign _14668_ = \bapg_rd.w_ptr_r [3] ? _14667_ : _14660_;
  assign _14669_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [13] : \MSYNC_1r1w.synth.nz.mem[304] [13];
  assign _14670_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [13] : \MSYNC_1r1w.synth.nz.mem[306] [13];
  assign _14671_ = \bapg_rd.w_ptr_r [1] ? _14670_ : _14669_;
  assign _14672_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [13] : \MSYNC_1r1w.synth.nz.mem[308] [13];
  assign _14673_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [13] : \MSYNC_1r1w.synth.nz.mem[310] [13];
  assign _14674_ = \bapg_rd.w_ptr_r [1] ? _14673_ : _14672_;
  assign _14675_ = \bapg_rd.w_ptr_r [2] ? _14674_ : _14671_;
  assign _14676_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [13] : \MSYNC_1r1w.synth.nz.mem[312] [13];
  assign _14677_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [13] : \MSYNC_1r1w.synth.nz.mem[314] [13];
  assign _14678_ = \bapg_rd.w_ptr_r [1] ? _14677_ : _14676_;
  assign _14679_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [13] : \MSYNC_1r1w.synth.nz.mem[316] [13];
  assign _14680_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [13] : \MSYNC_1r1w.synth.nz.mem[318] [13];
  assign _14681_ = \bapg_rd.w_ptr_r [1] ? _14680_ : _14679_;
  assign _14682_ = \bapg_rd.w_ptr_r [2] ? _14681_ : _14678_;
  assign _14683_ = \bapg_rd.w_ptr_r [3] ? _14682_ : _14675_;
  assign _14684_ = \bapg_rd.w_ptr_r [4] ? _14683_ : _14668_;
  assign _14685_ = \bapg_rd.w_ptr_r [5] ? _14684_ : _14653_;
  assign _14686_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [13] : \MSYNC_1r1w.synth.nz.mem[320] [13];
  assign _14687_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [13] : \MSYNC_1r1w.synth.nz.mem[322] [13];
  assign _14688_ = \bapg_rd.w_ptr_r [1] ? _14687_ : _14686_;
  assign _14689_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [13] : \MSYNC_1r1w.synth.nz.mem[324] [13];
  assign _14690_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [13] : \MSYNC_1r1w.synth.nz.mem[326] [13];
  assign _14691_ = \bapg_rd.w_ptr_r [1] ? _14690_ : _14689_;
  assign _14692_ = \bapg_rd.w_ptr_r [2] ? _14691_ : _14688_;
  assign _14693_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [13] : \MSYNC_1r1w.synth.nz.mem[328] [13];
  assign _14694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [13] : \MSYNC_1r1w.synth.nz.mem[330] [13];
  assign _14695_ = \bapg_rd.w_ptr_r [1] ? _14694_ : _14693_;
  assign _14696_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [13] : \MSYNC_1r1w.synth.nz.mem[332] [13];
  assign _14697_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [13] : \MSYNC_1r1w.synth.nz.mem[334] [13];
  assign _14698_ = \bapg_rd.w_ptr_r [1] ? _14697_ : _14696_;
  assign _14699_ = \bapg_rd.w_ptr_r [2] ? _14698_ : _14695_;
  assign _14700_ = \bapg_rd.w_ptr_r [3] ? _14699_ : _14692_;
  assign _14701_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [13] : \MSYNC_1r1w.synth.nz.mem[336] [13];
  assign _14702_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [13] : \MSYNC_1r1w.synth.nz.mem[338] [13];
  assign _14703_ = \bapg_rd.w_ptr_r [1] ? _14702_ : _14701_;
  assign _14704_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [13] : \MSYNC_1r1w.synth.nz.mem[340] [13];
  assign _14705_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [13] : \MSYNC_1r1w.synth.nz.mem[342] [13];
  assign _14706_ = \bapg_rd.w_ptr_r [1] ? _14705_ : _14704_;
  assign _14707_ = \bapg_rd.w_ptr_r [2] ? _14706_ : _14703_;
  assign _14708_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [13] : \MSYNC_1r1w.synth.nz.mem[344] [13];
  assign _14709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [13] : \MSYNC_1r1w.synth.nz.mem[346] [13];
  assign _14710_ = \bapg_rd.w_ptr_r [1] ? _14709_ : _14708_;
  assign _14711_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [13] : \MSYNC_1r1w.synth.nz.mem[348] [13];
  assign _14712_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [13] : \MSYNC_1r1w.synth.nz.mem[350] [13];
  assign _14713_ = \bapg_rd.w_ptr_r [1] ? _14712_ : _14711_;
  assign _14714_ = \bapg_rd.w_ptr_r [2] ? _14713_ : _14710_;
  assign _14715_ = \bapg_rd.w_ptr_r [3] ? _14714_ : _14707_;
  assign _14716_ = \bapg_rd.w_ptr_r [4] ? _14715_ : _14700_;
  assign _14717_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [13] : \MSYNC_1r1w.synth.nz.mem[352] [13];
  assign _14718_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [13] : \MSYNC_1r1w.synth.nz.mem[354] [13];
  assign _14719_ = \bapg_rd.w_ptr_r [1] ? _14718_ : _14717_;
  assign _14720_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [13] : \MSYNC_1r1w.synth.nz.mem[356] [13];
  assign _14721_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [13] : \MSYNC_1r1w.synth.nz.mem[358] [13];
  assign _14722_ = \bapg_rd.w_ptr_r [1] ? _14721_ : _14720_;
  assign _14723_ = \bapg_rd.w_ptr_r [2] ? _14722_ : _14719_;
  assign _14724_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [13] : \MSYNC_1r1w.synth.nz.mem[360] [13];
  assign _14725_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [13] : \MSYNC_1r1w.synth.nz.mem[362] [13];
  assign _14726_ = \bapg_rd.w_ptr_r [1] ? _14725_ : _14724_;
  assign _14727_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [13] : \MSYNC_1r1w.synth.nz.mem[364] [13];
  assign _14728_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [13] : \MSYNC_1r1w.synth.nz.mem[366] [13];
  assign _14729_ = \bapg_rd.w_ptr_r [1] ? _14728_ : _14727_;
  assign _14730_ = \bapg_rd.w_ptr_r [2] ? _14729_ : _14726_;
  assign _14731_ = \bapg_rd.w_ptr_r [3] ? _14730_ : _14723_;
  assign _14732_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [13] : \MSYNC_1r1w.synth.nz.mem[368] [13];
  assign _14733_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [13] : \MSYNC_1r1w.synth.nz.mem[370] [13];
  assign _14734_ = \bapg_rd.w_ptr_r [1] ? _14733_ : _14732_;
  assign _14735_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [13] : \MSYNC_1r1w.synth.nz.mem[372] [13];
  assign _14736_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [13] : \MSYNC_1r1w.synth.nz.mem[374] [13];
  assign _14737_ = \bapg_rd.w_ptr_r [1] ? _14736_ : _14735_;
  assign _14738_ = \bapg_rd.w_ptr_r [2] ? _14737_ : _14734_;
  assign _14739_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [13] : \MSYNC_1r1w.synth.nz.mem[376] [13];
  assign _14740_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [13] : \MSYNC_1r1w.synth.nz.mem[378] [13];
  assign _14741_ = \bapg_rd.w_ptr_r [1] ? _14740_ : _14739_;
  assign _14742_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [13] : \MSYNC_1r1w.synth.nz.mem[380] [13];
  assign _14743_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [13] : \MSYNC_1r1w.synth.nz.mem[382] [13];
  assign _14744_ = \bapg_rd.w_ptr_r [1] ? _14743_ : _14742_;
  assign _14745_ = \bapg_rd.w_ptr_r [2] ? _14744_ : _14741_;
  assign _14746_ = \bapg_rd.w_ptr_r [3] ? _14745_ : _14738_;
  assign _14747_ = \bapg_rd.w_ptr_r [4] ? _14746_ : _14731_;
  assign _14748_ = \bapg_rd.w_ptr_r [5] ? _14747_ : _14716_;
  assign _14749_ = \bapg_rd.w_ptr_r [6] ? _14748_ : _14685_;
  assign _14750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [13] : \MSYNC_1r1w.synth.nz.mem[384] [13];
  assign _14751_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [13] : \MSYNC_1r1w.synth.nz.mem[386] [13];
  assign _14752_ = \bapg_rd.w_ptr_r [1] ? _14751_ : _14750_;
  assign _14753_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [13] : \MSYNC_1r1w.synth.nz.mem[388] [13];
  assign _14754_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [13] : \MSYNC_1r1w.synth.nz.mem[390] [13];
  assign _14755_ = \bapg_rd.w_ptr_r [1] ? _14754_ : _14753_;
  assign _14756_ = \bapg_rd.w_ptr_r [2] ? _14755_ : _14752_;
  assign _14757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [13] : \MSYNC_1r1w.synth.nz.mem[392] [13];
  assign _14758_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [13] : \MSYNC_1r1w.synth.nz.mem[394] [13];
  assign _14759_ = \bapg_rd.w_ptr_r [1] ? _14758_ : _14757_;
  assign _14760_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [13] : \MSYNC_1r1w.synth.nz.mem[396] [13];
  assign _14761_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [13] : \MSYNC_1r1w.synth.nz.mem[398] [13];
  assign _14762_ = \bapg_rd.w_ptr_r [1] ? _14761_ : _14760_;
  assign _14763_ = \bapg_rd.w_ptr_r [2] ? _14762_ : _14759_;
  assign _14764_ = \bapg_rd.w_ptr_r [3] ? _14763_ : _14756_;
  assign _14765_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [13] : \MSYNC_1r1w.synth.nz.mem[400] [13];
  assign _14766_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [13] : \MSYNC_1r1w.synth.nz.mem[402] [13];
  assign _14767_ = \bapg_rd.w_ptr_r [1] ? _14766_ : _14765_;
  assign _14768_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [13] : \MSYNC_1r1w.synth.nz.mem[404] [13];
  assign _14769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [13] : \MSYNC_1r1w.synth.nz.mem[406] [13];
  assign _14770_ = \bapg_rd.w_ptr_r [1] ? _14769_ : _14768_;
  assign _14771_ = \bapg_rd.w_ptr_r [2] ? _14770_ : _14767_;
  assign _14772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [13] : \MSYNC_1r1w.synth.nz.mem[408] [13];
  assign _14773_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [13] : \MSYNC_1r1w.synth.nz.mem[410] [13];
  assign _14774_ = \bapg_rd.w_ptr_r [1] ? _14773_ : _14772_;
  assign _14775_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [13] : \MSYNC_1r1w.synth.nz.mem[412] [13];
  assign _14776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [13] : \MSYNC_1r1w.synth.nz.mem[414] [13];
  assign _14777_ = \bapg_rd.w_ptr_r [1] ? _14776_ : _14775_;
  assign _14778_ = \bapg_rd.w_ptr_r [2] ? _14777_ : _14774_;
  assign _14779_ = \bapg_rd.w_ptr_r [3] ? _14778_ : _14771_;
  assign _14780_ = \bapg_rd.w_ptr_r [4] ? _14779_ : _14764_;
  assign _14781_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [13] : \MSYNC_1r1w.synth.nz.mem[416] [13];
  assign _14782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [13] : \MSYNC_1r1w.synth.nz.mem[418] [13];
  assign _14783_ = \bapg_rd.w_ptr_r [1] ? _14782_ : _14781_;
  assign _14784_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [13] : \MSYNC_1r1w.synth.nz.mem[420] [13];
  assign _14785_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [13] : \MSYNC_1r1w.synth.nz.mem[422] [13];
  assign _14786_ = \bapg_rd.w_ptr_r [1] ? _14785_ : _14784_;
  assign _14787_ = \bapg_rd.w_ptr_r [2] ? _14786_ : _14783_;
  assign _14788_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [13] : \MSYNC_1r1w.synth.nz.mem[424] [13];
  assign _14789_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [13] : \MSYNC_1r1w.synth.nz.mem[426] [13];
  assign _14790_ = \bapg_rd.w_ptr_r [1] ? _14789_ : _14788_;
  assign _14791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [13] : \MSYNC_1r1w.synth.nz.mem[428] [13];
  assign _14792_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [13] : \MSYNC_1r1w.synth.nz.mem[430] [13];
  assign _14793_ = \bapg_rd.w_ptr_r [1] ? _14792_ : _14791_;
  assign _14794_ = \bapg_rd.w_ptr_r [2] ? _14793_ : _14790_;
  assign _14795_ = \bapg_rd.w_ptr_r [3] ? _14794_ : _14787_;
  assign _14796_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [13] : \MSYNC_1r1w.synth.nz.mem[432] [13];
  assign _14797_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [13] : \MSYNC_1r1w.synth.nz.mem[434] [13];
  assign _14798_ = \bapg_rd.w_ptr_r [1] ? _14797_ : _14796_;
  assign _14799_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [13] : \MSYNC_1r1w.synth.nz.mem[436] [13];
  assign _14800_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [13] : \MSYNC_1r1w.synth.nz.mem[438] [13];
  assign _14801_ = \bapg_rd.w_ptr_r [1] ? _14800_ : _14799_;
  assign _14802_ = \bapg_rd.w_ptr_r [2] ? _14801_ : _14798_;
  assign _14803_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [13] : \MSYNC_1r1w.synth.nz.mem[440] [13];
  assign _14804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [13] : \MSYNC_1r1w.synth.nz.mem[442] [13];
  assign _14805_ = \bapg_rd.w_ptr_r [1] ? _14804_ : _14803_;
  assign _14806_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [13] : \MSYNC_1r1w.synth.nz.mem[444] [13];
  assign _14807_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [13] : \MSYNC_1r1w.synth.nz.mem[446] [13];
  assign _14808_ = \bapg_rd.w_ptr_r [1] ? _14807_ : _14806_;
  assign _14809_ = \bapg_rd.w_ptr_r [2] ? _14808_ : _14805_;
  assign _14810_ = \bapg_rd.w_ptr_r [3] ? _14809_ : _14802_;
  assign _14811_ = \bapg_rd.w_ptr_r [4] ? _14810_ : _14795_;
  assign _14812_ = \bapg_rd.w_ptr_r [5] ? _14811_ : _14780_;
  assign _14813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [13] : \MSYNC_1r1w.synth.nz.mem[448] [13];
  assign _14814_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [13] : \MSYNC_1r1w.synth.nz.mem[450] [13];
  assign _14815_ = \bapg_rd.w_ptr_r [1] ? _14814_ : _14813_;
  assign _14816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [13] : \MSYNC_1r1w.synth.nz.mem[452] [13];
  assign _14817_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [13] : \MSYNC_1r1w.synth.nz.mem[454] [13];
  assign _14818_ = \bapg_rd.w_ptr_r [1] ? _14817_ : _14816_;
  assign _14819_ = \bapg_rd.w_ptr_r [2] ? _14818_ : _14815_;
  assign _14820_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [13] : \MSYNC_1r1w.synth.nz.mem[456] [13];
  assign _14821_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [13] : \MSYNC_1r1w.synth.nz.mem[458] [13];
  assign _14822_ = \bapg_rd.w_ptr_r [1] ? _14821_ : _14820_;
  assign _14823_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [13] : \MSYNC_1r1w.synth.nz.mem[460] [13];
  assign _14824_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [13] : \MSYNC_1r1w.synth.nz.mem[462] [13];
  assign _14825_ = \bapg_rd.w_ptr_r [1] ? _14824_ : _14823_;
  assign _14826_ = \bapg_rd.w_ptr_r [2] ? _14825_ : _14822_;
  assign _14827_ = \bapg_rd.w_ptr_r [3] ? _14826_ : _14819_;
  assign _14828_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [13] : \MSYNC_1r1w.synth.nz.mem[464] [13];
  assign _14829_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [13] : \MSYNC_1r1w.synth.nz.mem[466] [13];
  assign _14830_ = \bapg_rd.w_ptr_r [1] ? _14829_ : _14828_;
  assign _14831_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [13] : \MSYNC_1r1w.synth.nz.mem[468] [13];
  assign _14832_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [13] : \MSYNC_1r1w.synth.nz.mem[470] [13];
  assign _14833_ = \bapg_rd.w_ptr_r [1] ? _14832_ : _14831_;
  assign _14834_ = \bapg_rd.w_ptr_r [2] ? _14833_ : _14830_;
  assign _14835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [13] : \MSYNC_1r1w.synth.nz.mem[472] [13];
  assign _14836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [13] : \MSYNC_1r1w.synth.nz.mem[474] [13];
  assign _14837_ = \bapg_rd.w_ptr_r [1] ? _14836_ : _14835_;
  assign _14838_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [13] : \MSYNC_1r1w.synth.nz.mem[476] [13];
  assign _14839_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [13] : \MSYNC_1r1w.synth.nz.mem[478] [13];
  assign _14840_ = \bapg_rd.w_ptr_r [1] ? _14839_ : _14838_;
  assign _14841_ = \bapg_rd.w_ptr_r [2] ? _14840_ : _14837_;
  assign _14842_ = \bapg_rd.w_ptr_r [3] ? _14841_ : _14834_;
  assign _14843_ = \bapg_rd.w_ptr_r [4] ? _14842_ : _14827_;
  assign _14844_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [13] : \MSYNC_1r1w.synth.nz.mem[480] [13];
  assign _14845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [13] : \MSYNC_1r1w.synth.nz.mem[482] [13];
  assign _14846_ = \bapg_rd.w_ptr_r [1] ? _14845_ : _14844_;
  assign _14847_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [13] : \MSYNC_1r1w.synth.nz.mem[484] [13];
  assign _14848_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [13] : \MSYNC_1r1w.synth.nz.mem[486] [13];
  assign _14849_ = \bapg_rd.w_ptr_r [1] ? _14848_ : _14847_;
  assign _14850_ = \bapg_rd.w_ptr_r [2] ? _14849_ : _14846_;
  assign _14851_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [13] : \MSYNC_1r1w.synth.nz.mem[488] [13];
  assign _14852_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [13] : \MSYNC_1r1w.synth.nz.mem[490] [13];
  assign _14853_ = \bapg_rd.w_ptr_r [1] ? _14852_ : _14851_;
  assign _14854_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [13] : \MSYNC_1r1w.synth.nz.mem[492] [13];
  assign _14855_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [13] : \MSYNC_1r1w.synth.nz.mem[494] [13];
  assign _14856_ = \bapg_rd.w_ptr_r [1] ? _14855_ : _14854_;
  assign _14857_ = \bapg_rd.w_ptr_r [2] ? _14856_ : _14853_;
  assign _14858_ = \bapg_rd.w_ptr_r [3] ? _14857_ : _14850_;
  assign _14859_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [13] : \MSYNC_1r1w.synth.nz.mem[496] [13];
  assign _14860_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [13] : \MSYNC_1r1w.synth.nz.mem[498] [13];
  assign _14861_ = \bapg_rd.w_ptr_r [1] ? _14860_ : _14859_;
  assign _14862_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [13] : \MSYNC_1r1w.synth.nz.mem[500] [13];
  assign _14863_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [13] : \MSYNC_1r1w.synth.nz.mem[502] [13];
  assign _14864_ = \bapg_rd.w_ptr_r [1] ? _14863_ : _14862_;
  assign _14865_ = \bapg_rd.w_ptr_r [2] ? _14864_ : _14861_;
  assign _14866_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [13] : \MSYNC_1r1w.synth.nz.mem[504] [13];
  assign _14867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [13] : \MSYNC_1r1w.synth.nz.mem[506] [13];
  assign _14868_ = \bapg_rd.w_ptr_r [1] ? _14867_ : _14866_;
  assign _14869_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [13] : \MSYNC_1r1w.synth.nz.mem[508] [13];
  assign _14870_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [13] : \MSYNC_1r1w.synth.nz.mem[510] [13];
  assign _14871_ = \bapg_rd.w_ptr_r [1] ? _14870_ : _14869_;
  assign _14872_ = \bapg_rd.w_ptr_r [2] ? _14871_ : _14868_;
  assign _14873_ = \bapg_rd.w_ptr_r [3] ? _14872_ : _14865_;
  assign _14874_ = \bapg_rd.w_ptr_r [4] ? _14873_ : _14858_;
  assign _14875_ = \bapg_rd.w_ptr_r [5] ? _14874_ : _14843_;
  assign _14876_ = \bapg_rd.w_ptr_r [6] ? _14875_ : _14812_;
  assign _14877_ = \bapg_rd.w_ptr_r [7] ? _14876_ : _14749_;
  assign _14878_ = \bapg_rd.w_ptr_r [8] ? _14877_ : _14622_;
  assign _14879_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [13] : \MSYNC_1r1w.synth.nz.mem[512] [13];
  assign _14880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [13] : \MSYNC_1r1w.synth.nz.mem[514] [13];
  assign _14881_ = \bapg_rd.w_ptr_r [1] ? _14880_ : _14879_;
  assign _14882_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [13] : \MSYNC_1r1w.synth.nz.mem[516] [13];
  assign _14883_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [13] : \MSYNC_1r1w.synth.nz.mem[518] [13];
  assign _14884_ = \bapg_rd.w_ptr_r [1] ? _14883_ : _14882_;
  assign _14885_ = \bapg_rd.w_ptr_r [2] ? _14884_ : _14881_;
  assign _14886_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [13] : \MSYNC_1r1w.synth.nz.mem[520] [13];
  assign _14887_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [13] : \MSYNC_1r1w.synth.nz.mem[522] [13];
  assign _14888_ = \bapg_rd.w_ptr_r [1] ? _14887_ : _14886_;
  assign _14889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [13] : \MSYNC_1r1w.synth.nz.mem[524] [13];
  assign _14890_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [13] : \MSYNC_1r1w.synth.nz.mem[526] [13];
  assign _14891_ = \bapg_rd.w_ptr_r [1] ? _14890_ : _14889_;
  assign _14892_ = \bapg_rd.w_ptr_r [2] ? _14891_ : _14888_;
  assign _14893_ = \bapg_rd.w_ptr_r [3] ? _14892_ : _14885_;
  assign _14894_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [13] : \MSYNC_1r1w.synth.nz.mem[528] [13];
  assign _14895_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [13] : \MSYNC_1r1w.synth.nz.mem[530] [13];
  assign _14896_ = \bapg_rd.w_ptr_r [1] ? _14895_ : _14894_;
  assign _14897_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [13] : \MSYNC_1r1w.synth.nz.mem[532] [13];
  assign _14898_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [13] : \MSYNC_1r1w.synth.nz.mem[534] [13];
  assign _14899_ = \bapg_rd.w_ptr_r [1] ? _14898_ : _14897_;
  assign _14900_ = \bapg_rd.w_ptr_r [2] ? _14899_ : _14896_;
  assign _14901_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [13] : \MSYNC_1r1w.synth.nz.mem[536] [13];
  assign _14902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [13] : \MSYNC_1r1w.synth.nz.mem[538] [13];
  assign _14903_ = \bapg_rd.w_ptr_r [1] ? _14902_ : _14901_;
  assign _14904_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [13] : \MSYNC_1r1w.synth.nz.mem[540] [13];
  assign _14905_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [13] : \MSYNC_1r1w.synth.nz.mem[542] [13];
  assign _14906_ = \bapg_rd.w_ptr_r [1] ? _14905_ : _14904_;
  assign _14907_ = \bapg_rd.w_ptr_r [2] ? _14906_ : _14903_;
  assign _14908_ = \bapg_rd.w_ptr_r [3] ? _14907_ : _14900_;
  assign _14909_ = \bapg_rd.w_ptr_r [4] ? _14908_ : _14893_;
  assign _14910_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [13] : \MSYNC_1r1w.synth.nz.mem[544] [13];
  assign _14911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [13] : \MSYNC_1r1w.synth.nz.mem[546] [13];
  assign _14912_ = \bapg_rd.w_ptr_r [1] ? _14911_ : _14910_;
  assign _14913_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [13] : \MSYNC_1r1w.synth.nz.mem[548] [13];
  assign _14914_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [13] : \MSYNC_1r1w.synth.nz.mem[550] [13];
  assign _14915_ = \bapg_rd.w_ptr_r [1] ? _14914_ : _14913_;
  assign _14916_ = \bapg_rd.w_ptr_r [2] ? _14915_ : _14912_;
  assign _14917_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [13] : \MSYNC_1r1w.synth.nz.mem[552] [13];
  assign _14918_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [13] : \MSYNC_1r1w.synth.nz.mem[554] [13];
  assign _14919_ = \bapg_rd.w_ptr_r [1] ? _14918_ : _14917_;
  assign _14920_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [13] : \MSYNC_1r1w.synth.nz.mem[556] [13];
  assign _14921_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [13] : \MSYNC_1r1w.synth.nz.mem[558] [13];
  assign _14922_ = \bapg_rd.w_ptr_r [1] ? _14921_ : _14920_;
  assign _14923_ = \bapg_rd.w_ptr_r [2] ? _14922_ : _14919_;
  assign _14924_ = \bapg_rd.w_ptr_r [3] ? _14923_ : _14916_;
  assign _14925_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [13] : \MSYNC_1r1w.synth.nz.mem[560] [13];
  assign _14926_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [13] : \MSYNC_1r1w.synth.nz.mem[562] [13];
  assign _14927_ = \bapg_rd.w_ptr_r [1] ? _14926_ : _14925_;
  assign _14928_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [13] : \MSYNC_1r1w.synth.nz.mem[564] [13];
  assign _14929_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [13] : \MSYNC_1r1w.synth.nz.mem[566] [13];
  assign _14930_ = \bapg_rd.w_ptr_r [1] ? _14929_ : _14928_;
  assign _14931_ = \bapg_rd.w_ptr_r [2] ? _14930_ : _14927_;
  assign _14932_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [13] : \MSYNC_1r1w.synth.nz.mem[568] [13];
  assign _14933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [13] : \MSYNC_1r1w.synth.nz.mem[570] [13];
  assign _14934_ = \bapg_rd.w_ptr_r [1] ? _14933_ : _14932_;
  assign _14935_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [13] : \MSYNC_1r1w.synth.nz.mem[572] [13];
  assign _14936_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [13] : \MSYNC_1r1w.synth.nz.mem[574] [13];
  assign _14937_ = \bapg_rd.w_ptr_r [1] ? _14936_ : _14935_;
  assign _14938_ = \bapg_rd.w_ptr_r [2] ? _14937_ : _14934_;
  assign _14939_ = \bapg_rd.w_ptr_r [3] ? _14938_ : _14931_;
  assign _14940_ = \bapg_rd.w_ptr_r [4] ? _14939_ : _14924_;
  assign _14941_ = \bapg_rd.w_ptr_r [5] ? _14940_ : _14909_;
  assign _14942_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [13] : \MSYNC_1r1w.synth.nz.mem[576] [13];
  assign _14943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [13] : \MSYNC_1r1w.synth.nz.mem[578] [13];
  assign _14944_ = \bapg_rd.w_ptr_r [1] ? _14943_ : _14942_;
  assign _14945_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [13] : \MSYNC_1r1w.synth.nz.mem[580] [13];
  assign _14946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [13] : \MSYNC_1r1w.synth.nz.mem[582] [13];
  assign _14947_ = \bapg_rd.w_ptr_r [1] ? _14946_ : _14945_;
  assign _14948_ = \bapg_rd.w_ptr_r [2] ? _14947_ : _14944_;
  assign _14949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [13] : \MSYNC_1r1w.synth.nz.mem[584] [13];
  assign _14950_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [13] : \MSYNC_1r1w.synth.nz.mem[586] [13];
  assign _14951_ = \bapg_rd.w_ptr_r [1] ? _14950_ : _14949_;
  assign _14952_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [13] : \MSYNC_1r1w.synth.nz.mem[588] [13];
  assign _14953_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [13] : \MSYNC_1r1w.synth.nz.mem[590] [13];
  assign _14954_ = \bapg_rd.w_ptr_r [1] ? _14953_ : _14952_;
  assign _14955_ = \bapg_rd.w_ptr_r [2] ? _14954_ : _14951_;
  assign _14956_ = \bapg_rd.w_ptr_r [3] ? _14955_ : _14948_;
  assign _14957_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [13] : \MSYNC_1r1w.synth.nz.mem[592] [13];
  assign _14958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [13] : \MSYNC_1r1w.synth.nz.mem[594] [13];
  assign _14959_ = \bapg_rd.w_ptr_r [1] ? _14958_ : _14957_;
  assign _14960_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [13] : \MSYNC_1r1w.synth.nz.mem[596] [13];
  assign _14961_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [13] : \MSYNC_1r1w.synth.nz.mem[598] [13];
  assign _14962_ = \bapg_rd.w_ptr_r [1] ? _14961_ : _14960_;
  assign _14963_ = \bapg_rd.w_ptr_r [2] ? _14962_ : _14959_;
  assign _14964_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [13] : \MSYNC_1r1w.synth.nz.mem[600] [13];
  assign _14965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [13] : \MSYNC_1r1w.synth.nz.mem[602] [13];
  assign _14966_ = \bapg_rd.w_ptr_r [1] ? _14965_ : _14964_;
  assign _14967_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [13] : \MSYNC_1r1w.synth.nz.mem[604] [13];
  assign _14968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [13] : \MSYNC_1r1w.synth.nz.mem[606] [13];
  assign _14969_ = \bapg_rd.w_ptr_r [1] ? _14968_ : _14967_;
  assign _14970_ = \bapg_rd.w_ptr_r [2] ? _14969_ : _14966_;
  assign _14971_ = \bapg_rd.w_ptr_r [3] ? _14970_ : _14963_;
  assign _14972_ = \bapg_rd.w_ptr_r [4] ? _14971_ : _14956_;
  assign _14973_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [13] : \MSYNC_1r1w.synth.nz.mem[608] [13];
  assign _14974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [13] : \MSYNC_1r1w.synth.nz.mem[610] [13];
  assign _14975_ = \bapg_rd.w_ptr_r [1] ? _14974_ : _14973_;
  assign _14976_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [13] : \MSYNC_1r1w.synth.nz.mem[612] [13];
  assign _14977_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [13] : \MSYNC_1r1w.synth.nz.mem[614] [13];
  assign _14978_ = \bapg_rd.w_ptr_r [1] ? _14977_ : _14976_;
  assign _14979_ = \bapg_rd.w_ptr_r [2] ? _14978_ : _14975_;
  assign _14980_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [13] : \MSYNC_1r1w.synth.nz.mem[616] [13];
  assign _14981_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [13] : \MSYNC_1r1w.synth.nz.mem[618] [13];
  assign _14982_ = \bapg_rd.w_ptr_r [1] ? _14981_ : _14980_;
  assign _14983_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [13] : \MSYNC_1r1w.synth.nz.mem[620] [13];
  assign _14984_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [13] : \MSYNC_1r1w.synth.nz.mem[622] [13];
  assign _14985_ = \bapg_rd.w_ptr_r [1] ? _14984_ : _14983_;
  assign _14986_ = \bapg_rd.w_ptr_r [2] ? _14985_ : _14982_;
  assign _14987_ = \bapg_rd.w_ptr_r [3] ? _14986_ : _14979_;
  assign _14988_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [13] : \MSYNC_1r1w.synth.nz.mem[624] [13];
  assign _14989_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [13] : \MSYNC_1r1w.synth.nz.mem[626] [13];
  assign _14990_ = \bapg_rd.w_ptr_r [1] ? _14989_ : _14988_;
  assign _14991_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [13] : \MSYNC_1r1w.synth.nz.mem[628] [13];
  assign _14992_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [13] : \MSYNC_1r1w.synth.nz.mem[630] [13];
  assign _14993_ = \bapg_rd.w_ptr_r [1] ? _14992_ : _14991_;
  assign _14994_ = \bapg_rd.w_ptr_r [2] ? _14993_ : _14990_;
  assign _14995_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [13] : \MSYNC_1r1w.synth.nz.mem[632] [13];
  assign _14996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [13] : \MSYNC_1r1w.synth.nz.mem[634] [13];
  assign _14997_ = \bapg_rd.w_ptr_r [1] ? _14996_ : _14995_;
  assign _14998_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [13] : \MSYNC_1r1w.synth.nz.mem[636] [13];
  assign _14999_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [13] : \MSYNC_1r1w.synth.nz.mem[638] [13];
  assign _15000_ = \bapg_rd.w_ptr_r [1] ? _14999_ : _14998_;
  assign _15001_ = \bapg_rd.w_ptr_r [2] ? _15000_ : _14997_;
  assign _15002_ = \bapg_rd.w_ptr_r [3] ? _15001_ : _14994_;
  assign _15003_ = \bapg_rd.w_ptr_r [4] ? _15002_ : _14987_;
  assign _15004_ = \bapg_rd.w_ptr_r [5] ? _15003_ : _14972_;
  assign _15005_ = \bapg_rd.w_ptr_r [6] ? _15004_ : _14941_;
  assign _15006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [13] : \MSYNC_1r1w.synth.nz.mem[640] [13];
  assign _15007_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [13] : \MSYNC_1r1w.synth.nz.mem[642] [13];
  assign _15008_ = \bapg_rd.w_ptr_r [1] ? _15007_ : _15006_;
  assign _15009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [13] : \MSYNC_1r1w.synth.nz.mem[644] [13];
  assign _15010_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [13] : \MSYNC_1r1w.synth.nz.mem[646] [13];
  assign _15011_ = \bapg_rd.w_ptr_r [1] ? _15010_ : _15009_;
  assign _15012_ = \bapg_rd.w_ptr_r [2] ? _15011_ : _15008_;
  assign _15013_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [13] : \MSYNC_1r1w.synth.nz.mem[648] [13];
  assign _15014_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [13] : \MSYNC_1r1w.synth.nz.mem[650] [13];
  assign _15015_ = \bapg_rd.w_ptr_r [1] ? _15014_ : _15013_;
  assign _15016_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [13] : \MSYNC_1r1w.synth.nz.mem[652] [13];
  assign _15017_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [13] : \MSYNC_1r1w.synth.nz.mem[654] [13];
  assign _15018_ = \bapg_rd.w_ptr_r [1] ? _15017_ : _15016_;
  assign _15019_ = \bapg_rd.w_ptr_r [2] ? _15018_ : _15015_;
  assign _15020_ = \bapg_rd.w_ptr_r [3] ? _15019_ : _15012_;
  assign _15021_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [13] : \MSYNC_1r1w.synth.nz.mem[656] [13];
  assign _15022_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [13] : \MSYNC_1r1w.synth.nz.mem[658] [13];
  assign _15023_ = \bapg_rd.w_ptr_r [1] ? _15022_ : _15021_;
  assign _15024_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [13] : \MSYNC_1r1w.synth.nz.mem[660] [13];
  assign _15025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [13] : \MSYNC_1r1w.synth.nz.mem[662] [13];
  assign _15026_ = \bapg_rd.w_ptr_r [1] ? _15025_ : _15024_;
  assign _15027_ = \bapg_rd.w_ptr_r [2] ? _15026_ : _15023_;
  assign _15028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [13] : \MSYNC_1r1w.synth.nz.mem[664] [13];
  assign _15029_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [13] : \MSYNC_1r1w.synth.nz.mem[666] [13];
  assign _15030_ = \bapg_rd.w_ptr_r [1] ? _15029_ : _15028_;
  assign _15031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [13] : \MSYNC_1r1w.synth.nz.mem[668] [13];
  assign _15032_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [13] : \MSYNC_1r1w.synth.nz.mem[670] [13];
  assign _15033_ = \bapg_rd.w_ptr_r [1] ? _15032_ : _15031_;
  assign _15034_ = \bapg_rd.w_ptr_r [2] ? _15033_ : _15030_;
  assign _15035_ = \bapg_rd.w_ptr_r [3] ? _15034_ : _15027_;
  assign _15036_ = \bapg_rd.w_ptr_r [4] ? _15035_ : _15020_;
  assign _15037_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [13] : \MSYNC_1r1w.synth.nz.mem[672] [13];
  assign _15038_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [13] : \MSYNC_1r1w.synth.nz.mem[674] [13];
  assign _15039_ = \bapg_rd.w_ptr_r [1] ? _15038_ : _15037_;
  assign _15040_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [13] : \MSYNC_1r1w.synth.nz.mem[676] [13];
  assign _15041_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [13] : \MSYNC_1r1w.synth.nz.mem[678] [13];
  assign _15042_ = \bapg_rd.w_ptr_r [1] ? _15041_ : _15040_;
  assign _15043_ = \bapg_rd.w_ptr_r [2] ? _15042_ : _15039_;
  assign _15044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [13] : \MSYNC_1r1w.synth.nz.mem[680] [13];
  assign _15045_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [13] : \MSYNC_1r1w.synth.nz.mem[682] [13];
  assign _15046_ = \bapg_rd.w_ptr_r [1] ? _15045_ : _15044_;
  assign _15047_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [13] : \MSYNC_1r1w.synth.nz.mem[684] [13];
  assign _15048_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [13] : \MSYNC_1r1w.synth.nz.mem[686] [13];
  assign _15049_ = \bapg_rd.w_ptr_r [1] ? _15048_ : _15047_;
  assign _15050_ = \bapg_rd.w_ptr_r [2] ? _15049_ : _15046_;
  assign _15051_ = \bapg_rd.w_ptr_r [3] ? _15050_ : _15043_;
  assign _15052_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [13] : \MSYNC_1r1w.synth.nz.mem[688] [13];
  assign _15053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [13] : \MSYNC_1r1w.synth.nz.mem[690] [13];
  assign _15054_ = \bapg_rd.w_ptr_r [1] ? _15053_ : _15052_;
  assign _15055_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [13] : \MSYNC_1r1w.synth.nz.mem[692] [13];
  assign _15056_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [13] : \MSYNC_1r1w.synth.nz.mem[694] [13];
  assign _15057_ = \bapg_rd.w_ptr_r [1] ? _15056_ : _15055_;
  assign _15058_ = \bapg_rd.w_ptr_r [2] ? _15057_ : _15054_;
  assign _15059_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [13] : \MSYNC_1r1w.synth.nz.mem[696] [13];
  assign _15060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [13] : \MSYNC_1r1w.synth.nz.mem[698] [13];
  assign _15061_ = \bapg_rd.w_ptr_r [1] ? _15060_ : _15059_;
  assign _15062_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [13] : \MSYNC_1r1w.synth.nz.mem[700] [13];
  assign _15063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [13] : \MSYNC_1r1w.synth.nz.mem[702] [13];
  assign _15064_ = \bapg_rd.w_ptr_r [1] ? _15063_ : _15062_;
  assign _15065_ = \bapg_rd.w_ptr_r [2] ? _15064_ : _15061_;
  assign _15066_ = \bapg_rd.w_ptr_r [3] ? _15065_ : _15058_;
  assign _15067_ = \bapg_rd.w_ptr_r [4] ? _15066_ : _15051_;
  assign _15068_ = \bapg_rd.w_ptr_r [5] ? _15067_ : _15036_;
  assign _15069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [13] : \MSYNC_1r1w.synth.nz.mem[704] [13];
  assign _15070_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [13] : \MSYNC_1r1w.synth.nz.mem[706] [13];
  assign _15071_ = \bapg_rd.w_ptr_r [1] ? _15070_ : _15069_;
  assign _15072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [13] : \MSYNC_1r1w.synth.nz.mem[708] [13];
  assign _15073_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [13] : \MSYNC_1r1w.synth.nz.mem[710] [13];
  assign _15074_ = \bapg_rd.w_ptr_r [1] ? _15073_ : _15072_;
  assign _15075_ = \bapg_rd.w_ptr_r [2] ? _15074_ : _15071_;
  assign _15076_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [13] : \MSYNC_1r1w.synth.nz.mem[712] [13];
  assign _15077_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [13] : \MSYNC_1r1w.synth.nz.mem[714] [13];
  assign _15078_ = \bapg_rd.w_ptr_r [1] ? _15077_ : _15076_;
  assign _15079_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [13] : \MSYNC_1r1w.synth.nz.mem[716] [13];
  assign _15080_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [13] : \MSYNC_1r1w.synth.nz.mem[718] [13];
  assign _15081_ = \bapg_rd.w_ptr_r [1] ? _15080_ : _15079_;
  assign _15082_ = \bapg_rd.w_ptr_r [2] ? _15081_ : _15078_;
  assign _15083_ = \bapg_rd.w_ptr_r [3] ? _15082_ : _15075_;
  assign _15084_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [13] : \MSYNC_1r1w.synth.nz.mem[720] [13];
  assign _15085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [13] : \MSYNC_1r1w.synth.nz.mem[722] [13];
  assign _15086_ = \bapg_rd.w_ptr_r [1] ? _15085_ : _15084_;
  assign _15087_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [13] : \MSYNC_1r1w.synth.nz.mem[724] [13];
  assign _15088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [13] : \MSYNC_1r1w.synth.nz.mem[726] [13];
  assign _15089_ = \bapg_rd.w_ptr_r [1] ? _15088_ : _15087_;
  assign _15090_ = \bapg_rd.w_ptr_r [2] ? _15089_ : _15086_;
  assign _15091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [13] : \MSYNC_1r1w.synth.nz.mem[728] [13];
  assign _15092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [13] : \MSYNC_1r1w.synth.nz.mem[730] [13];
  assign _15093_ = \bapg_rd.w_ptr_r [1] ? _15092_ : _15091_;
  assign _15094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [13] : \MSYNC_1r1w.synth.nz.mem[732] [13];
  assign _15095_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [13] : \MSYNC_1r1w.synth.nz.mem[734] [13];
  assign _15096_ = \bapg_rd.w_ptr_r [1] ? _15095_ : _15094_;
  assign _15097_ = \bapg_rd.w_ptr_r [2] ? _15096_ : _15093_;
  assign _15098_ = \bapg_rd.w_ptr_r [3] ? _15097_ : _15090_;
  assign _15099_ = \bapg_rd.w_ptr_r [4] ? _15098_ : _15083_;
  assign _15100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [13] : \MSYNC_1r1w.synth.nz.mem[736] [13];
  assign _15101_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [13] : \MSYNC_1r1w.synth.nz.mem[738] [13];
  assign _15102_ = \bapg_rd.w_ptr_r [1] ? _15101_ : _15100_;
  assign _15103_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [13] : \MSYNC_1r1w.synth.nz.mem[740] [13];
  assign _15104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [13] : \MSYNC_1r1w.synth.nz.mem[742] [13];
  assign _15105_ = \bapg_rd.w_ptr_r [1] ? _15104_ : _15103_;
  assign _15106_ = \bapg_rd.w_ptr_r [2] ? _15105_ : _15102_;
  assign _15107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [13] : \MSYNC_1r1w.synth.nz.mem[744] [13];
  assign _15108_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [13] : \MSYNC_1r1w.synth.nz.mem[746] [13];
  assign _15109_ = \bapg_rd.w_ptr_r [1] ? _15108_ : _15107_;
  assign _15110_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [13] : \MSYNC_1r1w.synth.nz.mem[748] [13];
  assign _15111_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [13] : \MSYNC_1r1w.synth.nz.mem[750] [13];
  assign _15112_ = \bapg_rd.w_ptr_r [1] ? _15111_ : _15110_;
  assign _15113_ = \bapg_rd.w_ptr_r [2] ? _15112_ : _15109_;
  assign _15114_ = \bapg_rd.w_ptr_r [3] ? _15113_ : _15106_;
  assign _15115_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [13] : \MSYNC_1r1w.synth.nz.mem[752] [13];
  assign _15116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [13] : \MSYNC_1r1w.synth.nz.mem[754] [13];
  assign _15117_ = \bapg_rd.w_ptr_r [1] ? _15116_ : _15115_;
  assign _15118_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [13] : \MSYNC_1r1w.synth.nz.mem[756] [13];
  assign _15119_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [13] : \MSYNC_1r1w.synth.nz.mem[758] [13];
  assign _15120_ = \bapg_rd.w_ptr_r [1] ? _15119_ : _15118_;
  assign _15121_ = \bapg_rd.w_ptr_r [2] ? _15120_ : _15117_;
  assign _15122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [13] : \MSYNC_1r1w.synth.nz.mem[760] [13];
  assign _15123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [13] : \MSYNC_1r1w.synth.nz.mem[762] [13];
  assign _15124_ = \bapg_rd.w_ptr_r [1] ? _15123_ : _15122_;
  assign _15125_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [13] : \MSYNC_1r1w.synth.nz.mem[764] [13];
  assign _15126_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [13] : \MSYNC_1r1w.synth.nz.mem[766] [13];
  assign _15127_ = \bapg_rd.w_ptr_r [1] ? _15126_ : _15125_;
  assign _15128_ = \bapg_rd.w_ptr_r [2] ? _15127_ : _15124_;
  assign _15129_ = \bapg_rd.w_ptr_r [3] ? _15128_ : _15121_;
  assign _15130_ = \bapg_rd.w_ptr_r [4] ? _15129_ : _15114_;
  assign _15131_ = \bapg_rd.w_ptr_r [5] ? _15130_ : _15099_;
  assign _15132_ = \bapg_rd.w_ptr_r [6] ? _15131_ : _15068_;
  assign _15133_ = \bapg_rd.w_ptr_r [7] ? _15132_ : _15005_;
  assign _15134_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [13] : \MSYNC_1r1w.synth.nz.mem[768] [13];
  assign _15135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [13] : \MSYNC_1r1w.synth.nz.mem[770] [13];
  assign _15136_ = \bapg_rd.w_ptr_r [1] ? _15135_ : _15134_;
  assign _15137_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [13] : \MSYNC_1r1w.synth.nz.mem[772] [13];
  assign _15138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [13] : \MSYNC_1r1w.synth.nz.mem[774] [13];
  assign _15139_ = \bapg_rd.w_ptr_r [1] ? _15138_ : _15137_;
  assign _15140_ = \bapg_rd.w_ptr_r [2] ? _15139_ : _15136_;
  assign _15141_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [13] : \MSYNC_1r1w.synth.nz.mem[776] [13];
  assign _15142_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [13] : \MSYNC_1r1w.synth.nz.mem[778] [13];
  assign _15143_ = \bapg_rd.w_ptr_r [1] ? _15142_ : _15141_;
  assign _15144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [13] : \MSYNC_1r1w.synth.nz.mem[780] [13];
  assign _15145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [13] : \MSYNC_1r1w.synth.nz.mem[782] [13];
  assign _15146_ = \bapg_rd.w_ptr_r [1] ? _15145_ : _15144_;
  assign _15147_ = \bapg_rd.w_ptr_r [2] ? _15146_ : _15143_;
  assign _15148_ = \bapg_rd.w_ptr_r [3] ? _15147_ : _15140_;
  assign _15149_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [13] : \MSYNC_1r1w.synth.nz.mem[784] [13];
  assign _15150_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [13] : \MSYNC_1r1w.synth.nz.mem[786] [13];
  assign _15151_ = \bapg_rd.w_ptr_r [1] ? _15150_ : _15149_;
  assign _15152_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [13] : \MSYNC_1r1w.synth.nz.mem[788] [13];
  assign _15153_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [13] : \MSYNC_1r1w.synth.nz.mem[790] [13];
  assign _15154_ = \bapg_rd.w_ptr_r [1] ? _15153_ : _15152_;
  assign _15155_ = \bapg_rd.w_ptr_r [2] ? _15154_ : _15151_;
  assign _15156_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [13] : \MSYNC_1r1w.synth.nz.mem[792] [13];
  assign _15157_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [13] : \MSYNC_1r1w.synth.nz.mem[794] [13];
  assign _15158_ = \bapg_rd.w_ptr_r [1] ? _15157_ : _15156_;
  assign _15159_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [13] : \MSYNC_1r1w.synth.nz.mem[796] [13];
  assign _15160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [13] : \MSYNC_1r1w.synth.nz.mem[798] [13];
  assign _15161_ = \bapg_rd.w_ptr_r [1] ? _15160_ : _15159_;
  assign _15162_ = \bapg_rd.w_ptr_r [2] ? _15161_ : _15158_;
  assign _15163_ = \bapg_rd.w_ptr_r [3] ? _15162_ : _15155_;
  assign _15164_ = \bapg_rd.w_ptr_r [4] ? _15163_ : _15148_;
  assign _15165_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [13] : \MSYNC_1r1w.synth.nz.mem[800] [13];
  assign _15166_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [13] : \MSYNC_1r1w.synth.nz.mem[802] [13];
  assign _15167_ = \bapg_rd.w_ptr_r [1] ? _15166_ : _15165_;
  assign _15168_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [13] : \MSYNC_1r1w.synth.nz.mem[804] [13];
  assign _15169_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [13] : \MSYNC_1r1w.synth.nz.mem[806] [13];
  assign _15170_ = \bapg_rd.w_ptr_r [1] ? _15169_ : _15168_;
  assign _15171_ = \bapg_rd.w_ptr_r [2] ? _15170_ : _15167_;
  assign _15172_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [13] : \MSYNC_1r1w.synth.nz.mem[808] [13];
  assign _15173_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [13] : \MSYNC_1r1w.synth.nz.mem[810] [13];
  assign _15174_ = \bapg_rd.w_ptr_r [1] ? _15173_ : _15172_;
  assign _15175_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [13] : \MSYNC_1r1w.synth.nz.mem[812] [13];
  assign _15176_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [13] : \MSYNC_1r1w.synth.nz.mem[814] [13];
  assign _15177_ = \bapg_rd.w_ptr_r [1] ? _15176_ : _15175_;
  assign _15178_ = \bapg_rd.w_ptr_r [2] ? _15177_ : _15174_;
  assign _15179_ = \bapg_rd.w_ptr_r [3] ? _15178_ : _15171_;
  assign _15180_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [13] : \MSYNC_1r1w.synth.nz.mem[816] [13];
  assign _15181_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [13] : \MSYNC_1r1w.synth.nz.mem[818] [13];
  assign _15182_ = \bapg_rd.w_ptr_r [1] ? _15181_ : _15180_;
  assign _15183_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [13] : \MSYNC_1r1w.synth.nz.mem[820] [13];
  assign _15184_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [13] : \MSYNC_1r1w.synth.nz.mem[822] [13];
  assign _15185_ = \bapg_rd.w_ptr_r [1] ? _15184_ : _15183_;
  assign _15186_ = \bapg_rd.w_ptr_r [2] ? _15185_ : _15182_;
  assign _15187_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [13] : \MSYNC_1r1w.synth.nz.mem[824] [13];
  assign _15188_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [13] : \MSYNC_1r1w.synth.nz.mem[826] [13];
  assign _15189_ = \bapg_rd.w_ptr_r [1] ? _15188_ : _15187_;
  assign _15190_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [13] : \MSYNC_1r1w.synth.nz.mem[828] [13];
  assign _15191_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [13] : \MSYNC_1r1w.synth.nz.mem[830] [13];
  assign _15192_ = \bapg_rd.w_ptr_r [1] ? _15191_ : _15190_;
  assign _15193_ = \bapg_rd.w_ptr_r [2] ? _15192_ : _15189_;
  assign _15194_ = \bapg_rd.w_ptr_r [3] ? _15193_ : _15186_;
  assign _15195_ = \bapg_rd.w_ptr_r [4] ? _15194_ : _15179_;
  assign _15196_ = \bapg_rd.w_ptr_r [5] ? _15195_ : _15164_;
  assign _15197_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [13] : \MSYNC_1r1w.synth.nz.mem[832] [13];
  assign _15198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [13] : \MSYNC_1r1w.synth.nz.mem[834] [13];
  assign _15199_ = \bapg_rd.w_ptr_r [1] ? _15198_ : _15197_;
  assign _15200_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [13] : \MSYNC_1r1w.synth.nz.mem[836] [13];
  assign _15201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [13] : \MSYNC_1r1w.synth.nz.mem[838] [13];
  assign _15202_ = \bapg_rd.w_ptr_r [1] ? _15201_ : _15200_;
  assign _15203_ = \bapg_rd.w_ptr_r [2] ? _15202_ : _15199_;
  assign _15204_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [13] : \MSYNC_1r1w.synth.nz.mem[840] [13];
  assign _15205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [13] : \MSYNC_1r1w.synth.nz.mem[842] [13];
  assign _15206_ = \bapg_rd.w_ptr_r [1] ? _15205_ : _15204_;
  assign _15207_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [13] : \MSYNC_1r1w.synth.nz.mem[844] [13];
  assign _15208_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [13] : \MSYNC_1r1w.synth.nz.mem[846] [13];
  assign _15209_ = \bapg_rd.w_ptr_r [1] ? _15208_ : _15207_;
  assign _15210_ = \bapg_rd.w_ptr_r [2] ? _15209_ : _15206_;
  assign _15211_ = \bapg_rd.w_ptr_r [3] ? _15210_ : _15203_;
  assign _15212_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [13] : \MSYNC_1r1w.synth.nz.mem[848] [13];
  assign _15213_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [13] : \MSYNC_1r1w.synth.nz.mem[850] [13];
  assign _15214_ = \bapg_rd.w_ptr_r [1] ? _15213_ : _15212_;
  assign _15215_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [13] : \MSYNC_1r1w.synth.nz.mem[852] [13];
  assign _15216_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [13] : \MSYNC_1r1w.synth.nz.mem[854] [13];
  assign _15217_ = \bapg_rd.w_ptr_r [1] ? _15216_ : _15215_;
  assign _15218_ = \bapg_rd.w_ptr_r [2] ? _15217_ : _15214_;
  assign _15219_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [13] : \MSYNC_1r1w.synth.nz.mem[856] [13];
  assign _15220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [13] : \MSYNC_1r1w.synth.nz.mem[858] [13];
  assign _15221_ = \bapg_rd.w_ptr_r [1] ? _15220_ : _15219_;
  assign _15222_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [13] : \MSYNC_1r1w.synth.nz.mem[860] [13];
  assign _15223_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [13] : \MSYNC_1r1w.synth.nz.mem[862] [13];
  assign _15224_ = \bapg_rd.w_ptr_r [1] ? _15223_ : _15222_;
  assign _15225_ = \bapg_rd.w_ptr_r [2] ? _15224_ : _15221_;
  assign _15226_ = \bapg_rd.w_ptr_r [3] ? _15225_ : _15218_;
  assign _15227_ = \bapg_rd.w_ptr_r [4] ? _15226_ : _15211_;
  assign _15228_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [13] : \MSYNC_1r1w.synth.nz.mem[864] [13];
  assign _15229_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [13] : \MSYNC_1r1w.synth.nz.mem[866] [13];
  assign _15230_ = \bapg_rd.w_ptr_r [1] ? _15229_ : _15228_;
  assign _15231_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [13] : \MSYNC_1r1w.synth.nz.mem[868] [13];
  assign _15232_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [13] : \MSYNC_1r1w.synth.nz.mem[870] [13];
  assign _15233_ = \bapg_rd.w_ptr_r [1] ? _15232_ : _15231_;
  assign _15234_ = \bapg_rd.w_ptr_r [2] ? _15233_ : _15230_;
  assign _15235_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [13] : \MSYNC_1r1w.synth.nz.mem[872] [13];
  assign _15236_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [13] : \MSYNC_1r1w.synth.nz.mem[874] [13];
  assign _15237_ = \bapg_rd.w_ptr_r [1] ? _15236_ : _15235_;
  assign _15238_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [13] : \MSYNC_1r1w.synth.nz.mem[876] [13];
  assign _15239_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [13] : \MSYNC_1r1w.synth.nz.mem[878] [13];
  assign _15240_ = \bapg_rd.w_ptr_r [1] ? _15239_ : _15238_;
  assign _15241_ = \bapg_rd.w_ptr_r [2] ? _15240_ : _15237_;
  assign _15242_ = \bapg_rd.w_ptr_r [3] ? _15241_ : _15234_;
  assign _15243_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [13] : \MSYNC_1r1w.synth.nz.mem[880] [13];
  assign _15244_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [13] : \MSYNC_1r1w.synth.nz.mem[882] [13];
  assign _15245_ = \bapg_rd.w_ptr_r [1] ? _15244_ : _15243_;
  assign _15246_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [13] : \MSYNC_1r1w.synth.nz.mem[884] [13];
  assign _15247_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [13] : \MSYNC_1r1w.synth.nz.mem[886] [13];
  assign _15248_ = \bapg_rd.w_ptr_r [1] ? _15247_ : _15246_;
  assign _15249_ = \bapg_rd.w_ptr_r [2] ? _15248_ : _15245_;
  assign _15250_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [13] : \MSYNC_1r1w.synth.nz.mem[888] [13];
  assign _15251_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [13] : \MSYNC_1r1w.synth.nz.mem[890] [13];
  assign _15252_ = \bapg_rd.w_ptr_r [1] ? _15251_ : _15250_;
  assign _15253_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [13] : \MSYNC_1r1w.synth.nz.mem[892] [13];
  assign _15254_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [13] : \MSYNC_1r1w.synth.nz.mem[894] [13];
  assign _15255_ = \bapg_rd.w_ptr_r [1] ? _15254_ : _15253_;
  assign _15256_ = \bapg_rd.w_ptr_r [2] ? _15255_ : _15252_;
  assign _15257_ = \bapg_rd.w_ptr_r [3] ? _15256_ : _15249_;
  assign _15258_ = \bapg_rd.w_ptr_r [4] ? _15257_ : _15242_;
  assign _15259_ = \bapg_rd.w_ptr_r [5] ? _15258_ : _15227_;
  assign _15260_ = \bapg_rd.w_ptr_r [6] ? _15259_ : _15196_;
  assign _15261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [13] : \MSYNC_1r1w.synth.nz.mem[896] [13];
  assign _15262_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [13] : \MSYNC_1r1w.synth.nz.mem[898] [13];
  assign _15263_ = \bapg_rd.w_ptr_r [1] ? _15262_ : _15261_;
  assign _15264_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [13] : \MSYNC_1r1w.synth.nz.mem[900] [13];
  assign _15265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [13] : \MSYNC_1r1w.synth.nz.mem[902] [13];
  assign _15266_ = \bapg_rd.w_ptr_r [1] ? _15265_ : _15264_;
  assign _15267_ = \bapg_rd.w_ptr_r [2] ? _15266_ : _15263_;
  assign _15268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [13] : \MSYNC_1r1w.synth.nz.mem[904] [13];
  assign _15269_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [13] : \MSYNC_1r1w.synth.nz.mem[906] [13];
  assign _15270_ = \bapg_rd.w_ptr_r [1] ? _15269_ : _15268_;
  assign _15271_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [13] : \MSYNC_1r1w.synth.nz.mem[908] [13];
  assign _15272_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [13] : \MSYNC_1r1w.synth.nz.mem[910] [13];
  assign _15273_ = \bapg_rd.w_ptr_r [1] ? _15272_ : _15271_;
  assign _15274_ = \bapg_rd.w_ptr_r [2] ? _15273_ : _15270_;
  assign _15275_ = \bapg_rd.w_ptr_r [3] ? _15274_ : _15267_;
  assign _15276_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [13] : \MSYNC_1r1w.synth.nz.mem[912] [13];
  assign _15277_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [13] : \MSYNC_1r1w.synth.nz.mem[914] [13];
  assign _15278_ = \bapg_rd.w_ptr_r [1] ? _15277_ : _15276_;
  assign _15279_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [13] : \MSYNC_1r1w.synth.nz.mem[916] [13];
  assign _15280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [13] : \MSYNC_1r1w.synth.nz.mem[918] [13];
  assign _15281_ = \bapg_rd.w_ptr_r [1] ? _15280_ : _15279_;
  assign _15282_ = \bapg_rd.w_ptr_r [2] ? _15281_ : _15278_;
  assign _15283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [13] : \MSYNC_1r1w.synth.nz.mem[920] [13];
  assign _15284_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [13] : \MSYNC_1r1w.synth.nz.mem[922] [13];
  assign _15285_ = \bapg_rd.w_ptr_r [1] ? _15284_ : _15283_;
  assign _15286_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [13] : \MSYNC_1r1w.synth.nz.mem[924] [13];
  assign _15287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [13] : \MSYNC_1r1w.synth.nz.mem[926] [13];
  assign _15288_ = \bapg_rd.w_ptr_r [1] ? _15287_ : _15286_;
  assign _15289_ = \bapg_rd.w_ptr_r [2] ? _15288_ : _15285_;
  assign _15290_ = \bapg_rd.w_ptr_r [3] ? _15289_ : _15282_;
  assign _15291_ = \bapg_rd.w_ptr_r [4] ? _15290_ : _15275_;
  assign _15292_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [13] : \MSYNC_1r1w.synth.nz.mem[928] [13];
  assign _15293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [13] : \MSYNC_1r1w.synth.nz.mem[930] [13];
  assign _15294_ = \bapg_rd.w_ptr_r [1] ? _15293_ : _15292_;
  assign _15295_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [13] : \MSYNC_1r1w.synth.nz.mem[932] [13];
  assign _15296_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [13] : \MSYNC_1r1w.synth.nz.mem[934] [13];
  assign _15297_ = \bapg_rd.w_ptr_r [1] ? _15296_ : _15295_;
  assign _15298_ = \bapg_rd.w_ptr_r [2] ? _15297_ : _15294_;
  assign _15299_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [13] : \MSYNC_1r1w.synth.nz.mem[936] [13];
  assign _15300_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [13] : \MSYNC_1r1w.synth.nz.mem[938] [13];
  assign _15301_ = \bapg_rd.w_ptr_r [1] ? _15300_ : _15299_;
  assign _15302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [13] : \MSYNC_1r1w.synth.nz.mem[940] [13];
  assign _15303_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [13] : \MSYNC_1r1w.synth.nz.mem[942] [13];
  assign _15304_ = \bapg_rd.w_ptr_r [1] ? _15303_ : _15302_;
  assign _15305_ = \bapg_rd.w_ptr_r [2] ? _15304_ : _15301_;
  assign _15306_ = \bapg_rd.w_ptr_r [3] ? _15305_ : _15298_;
  assign _15307_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [13] : \MSYNC_1r1w.synth.nz.mem[944] [13];
  assign _15308_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [13] : \MSYNC_1r1w.synth.nz.mem[946] [13];
  assign _15309_ = \bapg_rd.w_ptr_r [1] ? _15308_ : _15307_;
  assign _15310_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [13] : \MSYNC_1r1w.synth.nz.mem[948] [13];
  assign _15311_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [13] : \MSYNC_1r1w.synth.nz.mem[950] [13];
  assign _15312_ = \bapg_rd.w_ptr_r [1] ? _15311_ : _15310_;
  assign _15313_ = \bapg_rd.w_ptr_r [2] ? _15312_ : _15309_;
  assign _15314_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [13] : \MSYNC_1r1w.synth.nz.mem[952] [13];
  assign _15315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [13] : \MSYNC_1r1w.synth.nz.mem[954] [13];
  assign _15316_ = \bapg_rd.w_ptr_r [1] ? _15315_ : _15314_;
  assign _15317_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [13] : \MSYNC_1r1w.synth.nz.mem[956] [13];
  assign _15318_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [13] : \MSYNC_1r1w.synth.nz.mem[958] [13];
  assign _15319_ = \bapg_rd.w_ptr_r [1] ? _15318_ : _15317_;
  assign _15320_ = \bapg_rd.w_ptr_r [2] ? _15319_ : _15316_;
  assign _15321_ = \bapg_rd.w_ptr_r [3] ? _15320_ : _15313_;
  assign _15322_ = \bapg_rd.w_ptr_r [4] ? _15321_ : _15306_;
  assign _15323_ = \bapg_rd.w_ptr_r [5] ? _15322_ : _15291_;
  assign _15324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [13] : \MSYNC_1r1w.synth.nz.mem[960] [13];
  assign _15325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [13] : \MSYNC_1r1w.synth.nz.mem[962] [13];
  assign _15326_ = \bapg_rd.w_ptr_r [1] ? _15325_ : _15324_;
  assign _15327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [13] : \MSYNC_1r1w.synth.nz.mem[964] [13];
  assign _15328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [13] : \MSYNC_1r1w.synth.nz.mem[966] [13];
  assign _15329_ = \bapg_rd.w_ptr_r [1] ? _15328_ : _15327_;
  assign _15330_ = \bapg_rd.w_ptr_r [2] ? _15329_ : _15326_;
  assign _15331_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [13] : \MSYNC_1r1w.synth.nz.mem[968] [13];
  assign _15332_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [13] : \MSYNC_1r1w.synth.nz.mem[970] [13];
  assign _15333_ = \bapg_rd.w_ptr_r [1] ? _15332_ : _15331_;
  assign _15334_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [13] : \MSYNC_1r1w.synth.nz.mem[972] [13];
  assign _15335_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [13] : \MSYNC_1r1w.synth.nz.mem[974] [13];
  assign _15336_ = \bapg_rd.w_ptr_r [1] ? _15335_ : _15334_;
  assign _15337_ = \bapg_rd.w_ptr_r [2] ? _15336_ : _15333_;
  assign _15338_ = \bapg_rd.w_ptr_r [3] ? _15337_ : _15330_;
  assign _15339_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [13] : \MSYNC_1r1w.synth.nz.mem[976] [13];
  assign _15340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [13] : \MSYNC_1r1w.synth.nz.mem[978] [13];
  assign _15341_ = \bapg_rd.w_ptr_r [1] ? _15340_ : _15339_;
  assign _15342_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [13] : \MSYNC_1r1w.synth.nz.mem[980] [13];
  assign _15343_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [13] : \MSYNC_1r1w.synth.nz.mem[982] [13];
  assign _15344_ = \bapg_rd.w_ptr_r [1] ? _15343_ : _15342_;
  assign _15345_ = \bapg_rd.w_ptr_r [2] ? _15344_ : _15341_;
  assign _15346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [13] : \MSYNC_1r1w.synth.nz.mem[984] [13];
  assign _15347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [13] : \MSYNC_1r1w.synth.nz.mem[986] [13];
  assign _15348_ = \bapg_rd.w_ptr_r [1] ? _15347_ : _15346_;
  assign _15349_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [13] : \MSYNC_1r1w.synth.nz.mem[988] [13];
  assign _15350_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [13] : \MSYNC_1r1w.synth.nz.mem[990] [13];
  assign _15351_ = \bapg_rd.w_ptr_r [1] ? _15350_ : _15349_;
  assign _15352_ = \bapg_rd.w_ptr_r [2] ? _15351_ : _15348_;
  assign _15353_ = \bapg_rd.w_ptr_r [3] ? _15352_ : _15345_;
  assign _15354_ = \bapg_rd.w_ptr_r [4] ? _15353_ : _15338_;
  assign _15355_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [13] : \MSYNC_1r1w.synth.nz.mem[992] [13];
  assign _15356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [13] : \MSYNC_1r1w.synth.nz.mem[994] [13];
  assign _15357_ = \bapg_rd.w_ptr_r [1] ? _15356_ : _15355_;
  assign _15358_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [13] : \MSYNC_1r1w.synth.nz.mem[996] [13];
  assign _15359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [13] : \MSYNC_1r1w.synth.nz.mem[998] [13];
  assign _15360_ = \bapg_rd.w_ptr_r [1] ? _15359_ : _15358_;
  assign _15361_ = \bapg_rd.w_ptr_r [2] ? _15360_ : _15357_;
  assign _15362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [13] : \MSYNC_1r1w.synth.nz.mem[1000] [13];
  assign _15363_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [13] : \MSYNC_1r1w.synth.nz.mem[1002] [13];
  assign _15364_ = \bapg_rd.w_ptr_r [1] ? _15363_ : _15362_;
  assign _15365_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [13] : \MSYNC_1r1w.synth.nz.mem[1004] [13];
  assign _15366_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [13] : \MSYNC_1r1w.synth.nz.mem[1006] [13];
  assign _15367_ = \bapg_rd.w_ptr_r [1] ? _15366_ : _15365_;
  assign _15368_ = \bapg_rd.w_ptr_r [2] ? _15367_ : _15364_;
  assign _15369_ = \bapg_rd.w_ptr_r [3] ? _15368_ : _15361_;
  assign _15370_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [13] : \MSYNC_1r1w.synth.nz.mem[1008] [13];
  assign _15371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [13] : \MSYNC_1r1w.synth.nz.mem[1010] [13];
  assign _15372_ = \bapg_rd.w_ptr_r [1] ? _15371_ : _15370_;
  assign _15373_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [13] : \MSYNC_1r1w.synth.nz.mem[1012] [13];
  assign _15374_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [13] : \MSYNC_1r1w.synth.nz.mem[1014] [13];
  assign _15375_ = \bapg_rd.w_ptr_r [1] ? _15374_ : _15373_;
  assign _15376_ = \bapg_rd.w_ptr_r [2] ? _15375_ : _15372_;
  assign _15377_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [13] : \MSYNC_1r1w.synth.nz.mem[1016] [13];
  assign _15378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [13] : \MSYNC_1r1w.synth.nz.mem[1018] [13];
  assign _15379_ = \bapg_rd.w_ptr_r [1] ? _15378_ : _15377_;
  assign _15380_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [13] : \MSYNC_1r1w.synth.nz.mem[1020] [13];
  assign _15381_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [13] : \MSYNC_1r1w.synth.nz.mem[1022] [13];
  assign _15382_ = \bapg_rd.w_ptr_r [1] ? _15381_ : _15380_;
  assign _15383_ = \bapg_rd.w_ptr_r [2] ? _15382_ : _15379_;
  assign _15384_ = \bapg_rd.w_ptr_r [3] ? _15383_ : _15376_;
  assign _15385_ = \bapg_rd.w_ptr_r [4] ? _15384_ : _15369_;
  assign _15386_ = \bapg_rd.w_ptr_r [5] ? _15385_ : _15354_;
  assign _15387_ = \bapg_rd.w_ptr_r [6] ? _15386_ : _15323_;
  assign _15388_ = \bapg_rd.w_ptr_r [7] ? _15387_ : _15260_;
  assign _15389_ = \bapg_rd.w_ptr_r [8] ? _15388_ : _15133_;
  assign r_data_o[13] = \bapg_rd.w_ptr_r [9] ? _15389_ : _14878_;
  assign _15390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [14] : \MSYNC_1r1w.synth.nz.mem[0] [14];
  assign _15391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [14] : \MSYNC_1r1w.synth.nz.mem[2] [14];
  assign _15392_ = \bapg_rd.w_ptr_r [1] ? _15391_ : _15390_;
  assign _15393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [14] : \MSYNC_1r1w.synth.nz.mem[4] [14];
  assign _15394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [14] : \MSYNC_1r1w.synth.nz.mem[6] [14];
  assign _15395_ = \bapg_rd.w_ptr_r [1] ? _15394_ : _15393_;
  assign _15396_ = \bapg_rd.w_ptr_r [2] ? _15395_ : _15392_;
  assign _15397_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [14] : \MSYNC_1r1w.synth.nz.mem[8] [14];
  assign _15398_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [14] : \MSYNC_1r1w.synth.nz.mem[10] [14];
  assign _15399_ = \bapg_rd.w_ptr_r [1] ? _15398_ : _15397_;
  assign _15400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [14] : \MSYNC_1r1w.synth.nz.mem[12] [14];
  assign _15401_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [14] : \MSYNC_1r1w.synth.nz.mem[14] [14];
  assign _15402_ = \bapg_rd.w_ptr_r [1] ? _15401_ : _15400_;
  assign _15403_ = \bapg_rd.w_ptr_r [2] ? _15402_ : _15399_;
  assign _15404_ = \bapg_rd.w_ptr_r [3] ? _15403_ : _15396_;
  assign _15405_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [14] : \MSYNC_1r1w.synth.nz.mem[16] [14];
  assign _15406_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [14] : \MSYNC_1r1w.synth.nz.mem[18] [14];
  assign _15407_ = \bapg_rd.w_ptr_r [1] ? _15406_ : _15405_;
  assign _15408_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [14] : \MSYNC_1r1w.synth.nz.mem[20] [14];
  assign _15409_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [14] : \MSYNC_1r1w.synth.nz.mem[22] [14];
  assign _15410_ = \bapg_rd.w_ptr_r [1] ? _15409_ : _15408_;
  assign _15411_ = \bapg_rd.w_ptr_r [2] ? _15410_ : _15407_;
  assign _15412_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [14] : \MSYNC_1r1w.synth.nz.mem[24] [14];
  assign _15413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [14] : \MSYNC_1r1w.synth.nz.mem[26] [14];
  assign _15414_ = \bapg_rd.w_ptr_r [1] ? _15413_ : _15412_;
  assign _15415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [14] : \MSYNC_1r1w.synth.nz.mem[28] [14];
  assign _15416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [14] : \MSYNC_1r1w.synth.nz.mem[30] [14];
  assign _15417_ = \bapg_rd.w_ptr_r [1] ? _15416_ : _15415_;
  assign _15418_ = \bapg_rd.w_ptr_r [2] ? _15417_ : _15414_;
  assign _15419_ = \bapg_rd.w_ptr_r [3] ? _15418_ : _15411_;
  assign _15420_ = \bapg_rd.w_ptr_r [4] ? _15419_ : _15404_;
  assign _15421_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [14] : \MSYNC_1r1w.synth.nz.mem[32] [14];
  assign _15422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [14] : \MSYNC_1r1w.synth.nz.mem[34] [14];
  assign _15423_ = \bapg_rd.w_ptr_r [1] ? _15422_ : _15421_;
  assign _15424_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [14] : \MSYNC_1r1w.synth.nz.mem[36] [14];
  assign _15425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [14] : \MSYNC_1r1w.synth.nz.mem[38] [14];
  assign _15426_ = \bapg_rd.w_ptr_r [1] ? _15425_ : _15424_;
  assign _15427_ = \bapg_rd.w_ptr_r [2] ? _15426_ : _15423_;
  assign _15428_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [14] : \MSYNC_1r1w.synth.nz.mem[40] [14];
  assign _15429_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [14] : \MSYNC_1r1w.synth.nz.mem[42] [14];
  assign _15430_ = \bapg_rd.w_ptr_r [1] ? _15429_ : _15428_;
  assign _15431_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [14] : \MSYNC_1r1w.synth.nz.mem[44] [14];
  assign _15432_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [14] : \MSYNC_1r1w.synth.nz.mem[46] [14];
  assign _15433_ = \bapg_rd.w_ptr_r [1] ? _15432_ : _15431_;
  assign _15434_ = \bapg_rd.w_ptr_r [2] ? _15433_ : _15430_;
  assign _15435_ = \bapg_rd.w_ptr_r [3] ? _15434_ : _15427_;
  assign _15436_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [14] : \MSYNC_1r1w.synth.nz.mem[48] [14];
  assign _15437_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [14] : \MSYNC_1r1w.synth.nz.mem[50] [14];
  assign _15438_ = \bapg_rd.w_ptr_r [1] ? _15437_ : _15436_;
  assign _15439_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [14] : \MSYNC_1r1w.synth.nz.mem[52] [14];
  assign _15440_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [14] : \MSYNC_1r1w.synth.nz.mem[54] [14];
  assign _15441_ = \bapg_rd.w_ptr_r [1] ? _15440_ : _15439_;
  assign _15442_ = \bapg_rd.w_ptr_r [2] ? _15441_ : _15438_;
  assign _15443_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [14] : \MSYNC_1r1w.synth.nz.mem[56] [14];
  assign _15444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [14] : \MSYNC_1r1w.synth.nz.mem[58] [14];
  assign _15445_ = \bapg_rd.w_ptr_r [1] ? _15444_ : _15443_;
  assign _15446_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [14] : \MSYNC_1r1w.synth.nz.mem[60] [14];
  assign _15447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [14] : \MSYNC_1r1w.synth.nz.mem[62] [14];
  assign _15448_ = \bapg_rd.w_ptr_r [1] ? _15447_ : _15446_;
  assign _15449_ = \bapg_rd.w_ptr_r [2] ? _15448_ : _15445_;
  assign _15450_ = \bapg_rd.w_ptr_r [3] ? _15449_ : _15442_;
  assign _15451_ = \bapg_rd.w_ptr_r [4] ? _15450_ : _15435_;
  assign _15452_ = \bapg_rd.w_ptr_r [5] ? _15451_ : _15420_;
  assign _15453_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [14] : \MSYNC_1r1w.synth.nz.mem[64] [14];
  assign _15454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [14] : \MSYNC_1r1w.synth.nz.mem[66] [14];
  assign _15455_ = \bapg_rd.w_ptr_r [1] ? _15454_ : _15453_;
  assign _15456_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [14] : \MSYNC_1r1w.synth.nz.mem[68] [14];
  assign _15457_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [14] : \MSYNC_1r1w.synth.nz.mem[70] [14];
  assign _15458_ = \bapg_rd.w_ptr_r [1] ? _15457_ : _15456_;
  assign _15459_ = \bapg_rd.w_ptr_r [2] ? _15458_ : _15455_;
  assign _15460_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [14] : \MSYNC_1r1w.synth.nz.mem[72] [14];
  assign _15461_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [14] : \MSYNC_1r1w.synth.nz.mem[74] [14];
  assign _15462_ = \bapg_rd.w_ptr_r [1] ? _15461_ : _15460_;
  assign _15463_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [14] : \MSYNC_1r1w.synth.nz.mem[76] [14];
  assign _15464_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [14] : \MSYNC_1r1w.synth.nz.mem[78] [14];
  assign _15465_ = \bapg_rd.w_ptr_r [1] ? _15464_ : _15463_;
  assign _15466_ = \bapg_rd.w_ptr_r [2] ? _15465_ : _15462_;
  assign _15467_ = \bapg_rd.w_ptr_r [3] ? _15466_ : _15459_;
  assign _15468_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [14] : \MSYNC_1r1w.synth.nz.mem[80] [14];
  assign _15469_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [14] : \MSYNC_1r1w.synth.nz.mem[82] [14];
  assign _15470_ = \bapg_rd.w_ptr_r [1] ? _15469_ : _15468_;
  assign _15471_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [14] : \MSYNC_1r1w.synth.nz.mem[84] [14];
  assign _15472_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [14] : \MSYNC_1r1w.synth.nz.mem[86] [14];
  assign _15473_ = \bapg_rd.w_ptr_r [1] ? _15472_ : _15471_;
  assign _15474_ = \bapg_rd.w_ptr_r [2] ? _15473_ : _15470_;
  assign _15475_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [14] : \MSYNC_1r1w.synth.nz.mem[88] [14];
  assign _15476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [14] : \MSYNC_1r1w.synth.nz.mem[90] [14];
  assign _15477_ = \bapg_rd.w_ptr_r [1] ? _15476_ : _15475_;
  assign _15478_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [14] : \MSYNC_1r1w.synth.nz.mem[92] [14];
  assign _15479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [14] : \MSYNC_1r1w.synth.nz.mem[94] [14];
  assign _15480_ = \bapg_rd.w_ptr_r [1] ? _15479_ : _15478_;
  assign _15481_ = \bapg_rd.w_ptr_r [2] ? _15480_ : _15477_;
  assign _15482_ = \bapg_rd.w_ptr_r [3] ? _15481_ : _15474_;
  assign _15483_ = \bapg_rd.w_ptr_r [4] ? _15482_ : _15467_;
  assign _15484_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [14] : \MSYNC_1r1w.synth.nz.mem[96] [14];
  assign _15485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [14] : \MSYNC_1r1w.synth.nz.mem[98] [14];
  assign _15486_ = \bapg_rd.w_ptr_r [1] ? _15485_ : _15484_;
  assign _15487_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [14] : \MSYNC_1r1w.synth.nz.mem[100] [14];
  assign _15488_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [14] : \MSYNC_1r1w.synth.nz.mem[102] [14];
  assign _15489_ = \bapg_rd.w_ptr_r [1] ? _15488_ : _15487_;
  assign _15490_ = \bapg_rd.w_ptr_r [2] ? _15489_ : _15486_;
  assign _15491_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [14] : \MSYNC_1r1w.synth.nz.mem[104] [14];
  assign _15492_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [14] : \MSYNC_1r1w.synth.nz.mem[106] [14];
  assign _15493_ = \bapg_rd.w_ptr_r [1] ? _15492_ : _15491_;
  assign _15494_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [14] : \MSYNC_1r1w.synth.nz.mem[108] [14];
  assign _15495_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [14] : \MSYNC_1r1w.synth.nz.mem[110] [14];
  assign _15496_ = \bapg_rd.w_ptr_r [1] ? _15495_ : _15494_;
  assign _15497_ = \bapg_rd.w_ptr_r [2] ? _15496_ : _15493_;
  assign _15498_ = \bapg_rd.w_ptr_r [3] ? _15497_ : _15490_;
  assign _15499_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [14] : \MSYNC_1r1w.synth.nz.mem[112] [14];
  assign _15500_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [14] : \MSYNC_1r1w.synth.nz.mem[114] [14];
  assign _15501_ = \bapg_rd.w_ptr_r [1] ? _15500_ : _15499_;
  assign _15502_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [14] : \MSYNC_1r1w.synth.nz.mem[116] [14];
  assign _15503_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [14] : \MSYNC_1r1w.synth.nz.mem[118] [14];
  assign _15504_ = \bapg_rd.w_ptr_r [1] ? _15503_ : _15502_;
  assign _15505_ = \bapg_rd.w_ptr_r [2] ? _15504_ : _15501_;
  assign _15506_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [14] : \MSYNC_1r1w.synth.nz.mem[120] [14];
  assign _15507_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [14] : \MSYNC_1r1w.synth.nz.mem[122] [14];
  assign _15508_ = \bapg_rd.w_ptr_r [1] ? _15507_ : _15506_;
  assign _15509_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [14] : \MSYNC_1r1w.synth.nz.mem[124] [14];
  assign _15510_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [14] : \MSYNC_1r1w.synth.nz.mem[126] [14];
  assign _15511_ = \bapg_rd.w_ptr_r [1] ? _15510_ : _15509_;
  assign _15512_ = \bapg_rd.w_ptr_r [2] ? _15511_ : _15508_;
  assign _15513_ = \bapg_rd.w_ptr_r [3] ? _15512_ : _15505_;
  assign _15514_ = \bapg_rd.w_ptr_r [4] ? _15513_ : _15498_;
  assign _15515_ = \bapg_rd.w_ptr_r [5] ? _15514_ : _15483_;
  assign _15516_ = \bapg_rd.w_ptr_r [6] ? _15515_ : _15452_;
  assign _15517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [14] : \MSYNC_1r1w.synth.nz.mem[128] [14];
  assign _15518_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [14] : \MSYNC_1r1w.synth.nz.mem[130] [14];
  assign _15519_ = \bapg_rd.w_ptr_r [1] ? _15518_ : _15517_;
  assign _15520_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [14] : \MSYNC_1r1w.synth.nz.mem[132] [14];
  assign _15521_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [14] : \MSYNC_1r1w.synth.nz.mem[134] [14];
  assign _15522_ = \bapg_rd.w_ptr_r [1] ? _15521_ : _15520_;
  assign _15523_ = \bapg_rd.w_ptr_r [2] ? _15522_ : _15519_;
  assign _15524_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [14] : \MSYNC_1r1w.synth.nz.mem[136] [14];
  assign _15525_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [14] : \MSYNC_1r1w.synth.nz.mem[138] [14];
  assign _15526_ = \bapg_rd.w_ptr_r [1] ? _15525_ : _15524_;
  assign _15527_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [14] : \MSYNC_1r1w.synth.nz.mem[140] [14];
  assign _15528_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [14] : \MSYNC_1r1w.synth.nz.mem[142] [14];
  assign _15529_ = \bapg_rd.w_ptr_r [1] ? _15528_ : _15527_;
  assign _15530_ = \bapg_rd.w_ptr_r [2] ? _15529_ : _15526_;
  assign _15531_ = \bapg_rd.w_ptr_r [3] ? _15530_ : _15523_;
  assign _15532_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [14] : \MSYNC_1r1w.synth.nz.mem[144] [14];
  assign _15533_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [14] : \MSYNC_1r1w.synth.nz.mem[146] [14];
  assign _15534_ = \bapg_rd.w_ptr_r [1] ? _15533_ : _15532_;
  assign _15535_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [14] : \MSYNC_1r1w.synth.nz.mem[148] [14];
  assign _15536_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [14] : \MSYNC_1r1w.synth.nz.mem[150] [14];
  assign _15537_ = \bapg_rd.w_ptr_r [1] ? _15536_ : _15535_;
  assign _15538_ = \bapg_rd.w_ptr_r [2] ? _15537_ : _15534_;
  assign _15539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [14] : \MSYNC_1r1w.synth.nz.mem[152] [14];
  assign _15540_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [14] : \MSYNC_1r1w.synth.nz.mem[154] [14];
  assign _15541_ = \bapg_rd.w_ptr_r [1] ? _15540_ : _15539_;
  assign _15542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [14] : \MSYNC_1r1w.synth.nz.mem[156] [14];
  assign _15543_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [14] : \MSYNC_1r1w.synth.nz.mem[158] [14];
  assign _15544_ = \bapg_rd.w_ptr_r [1] ? _15543_ : _15542_;
  assign _15545_ = \bapg_rd.w_ptr_r [2] ? _15544_ : _15541_;
  assign _15546_ = \bapg_rd.w_ptr_r [3] ? _15545_ : _15538_;
  assign _15547_ = \bapg_rd.w_ptr_r [4] ? _15546_ : _15531_;
  assign _15548_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [14] : \MSYNC_1r1w.synth.nz.mem[160] [14];
  assign _15549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [14] : \MSYNC_1r1w.synth.nz.mem[162] [14];
  assign _15550_ = \bapg_rd.w_ptr_r [1] ? _15549_ : _15548_;
  assign _15551_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [14] : \MSYNC_1r1w.synth.nz.mem[164] [14];
  assign _15552_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [14] : \MSYNC_1r1w.synth.nz.mem[166] [14];
  assign _15553_ = \bapg_rd.w_ptr_r [1] ? _15552_ : _15551_;
  assign _15554_ = \bapg_rd.w_ptr_r [2] ? _15553_ : _15550_;
  assign _15555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [14] : \MSYNC_1r1w.synth.nz.mem[168] [14];
  assign _15556_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [14] : \MSYNC_1r1w.synth.nz.mem[170] [14];
  assign _15557_ = \bapg_rd.w_ptr_r [1] ? _15556_ : _15555_;
  assign _15558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [14] : \MSYNC_1r1w.synth.nz.mem[172] [14];
  assign _15559_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [14] : \MSYNC_1r1w.synth.nz.mem[174] [14];
  assign _15560_ = \bapg_rd.w_ptr_r [1] ? _15559_ : _15558_;
  assign _15561_ = \bapg_rd.w_ptr_r [2] ? _15560_ : _15557_;
  assign _15562_ = \bapg_rd.w_ptr_r [3] ? _15561_ : _15554_;
  assign _15563_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [14] : \MSYNC_1r1w.synth.nz.mem[176] [14];
  assign _15564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [14] : \MSYNC_1r1w.synth.nz.mem[178] [14];
  assign _15565_ = \bapg_rd.w_ptr_r [1] ? _15564_ : _15563_;
  assign _15566_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [14] : \MSYNC_1r1w.synth.nz.mem[180] [14];
  assign _15567_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [14] : \MSYNC_1r1w.synth.nz.mem[182] [14];
  assign _15568_ = \bapg_rd.w_ptr_r [1] ? _15567_ : _15566_;
  assign _15569_ = \bapg_rd.w_ptr_r [2] ? _15568_ : _15565_;
  assign _15570_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [14] : \MSYNC_1r1w.synth.nz.mem[184] [14];
  assign _15571_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [14] : \MSYNC_1r1w.synth.nz.mem[186] [14];
  assign _15572_ = \bapg_rd.w_ptr_r [1] ? _15571_ : _15570_;
  assign _15573_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [14] : \MSYNC_1r1w.synth.nz.mem[188] [14];
  assign _15574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [14] : \MSYNC_1r1w.synth.nz.mem[190] [14];
  assign _15575_ = \bapg_rd.w_ptr_r [1] ? _15574_ : _15573_;
  assign _15576_ = \bapg_rd.w_ptr_r [2] ? _15575_ : _15572_;
  assign _15577_ = \bapg_rd.w_ptr_r [3] ? _15576_ : _15569_;
  assign _15578_ = \bapg_rd.w_ptr_r [4] ? _15577_ : _15562_;
  assign _15579_ = \bapg_rd.w_ptr_r [5] ? _15578_ : _15547_;
  assign _15580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [14] : \MSYNC_1r1w.synth.nz.mem[192] [14];
  assign _15581_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [14] : \MSYNC_1r1w.synth.nz.mem[194] [14];
  assign _15582_ = \bapg_rd.w_ptr_r [1] ? _15581_ : _15580_;
  assign _15583_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [14] : \MSYNC_1r1w.synth.nz.mem[196] [14];
  assign _15584_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [14] : \MSYNC_1r1w.synth.nz.mem[198] [14];
  assign _15585_ = \bapg_rd.w_ptr_r [1] ? _15584_ : _15583_;
  assign _15586_ = \bapg_rd.w_ptr_r [2] ? _15585_ : _15582_;
  assign _15587_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [14] : \MSYNC_1r1w.synth.nz.mem[200] [14];
  assign _15588_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [14] : \MSYNC_1r1w.synth.nz.mem[202] [14];
  assign _15589_ = \bapg_rd.w_ptr_r [1] ? _15588_ : _15587_;
  assign _15590_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [14] : \MSYNC_1r1w.synth.nz.mem[204] [14];
  assign _15591_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [14] : \MSYNC_1r1w.synth.nz.mem[206] [14];
  assign _15592_ = \bapg_rd.w_ptr_r [1] ? _15591_ : _15590_;
  assign _15593_ = \bapg_rd.w_ptr_r [2] ? _15592_ : _15589_;
  assign _15594_ = \bapg_rd.w_ptr_r [3] ? _15593_ : _15586_;
  assign _15595_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [14] : \MSYNC_1r1w.synth.nz.mem[208] [14];
  assign _15596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [14] : \MSYNC_1r1w.synth.nz.mem[210] [14];
  assign _15597_ = \bapg_rd.w_ptr_r [1] ? _15596_ : _15595_;
  assign _15598_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [14] : \MSYNC_1r1w.synth.nz.mem[212] [14];
  assign _15599_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [14] : \MSYNC_1r1w.synth.nz.mem[214] [14];
  assign _15600_ = \bapg_rd.w_ptr_r [1] ? _15599_ : _15598_;
  assign _15601_ = \bapg_rd.w_ptr_r [2] ? _15600_ : _15597_;
  assign _15602_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [14] : \MSYNC_1r1w.synth.nz.mem[216] [14];
  assign _15603_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [14] : \MSYNC_1r1w.synth.nz.mem[218] [14];
  assign _15604_ = \bapg_rd.w_ptr_r [1] ? _15603_ : _15602_;
  assign _15605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [14] : \MSYNC_1r1w.synth.nz.mem[220] [14];
  assign _15606_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [14] : \MSYNC_1r1w.synth.nz.mem[222] [14];
  assign _15607_ = \bapg_rd.w_ptr_r [1] ? _15606_ : _15605_;
  assign _15608_ = \bapg_rd.w_ptr_r [2] ? _15607_ : _15604_;
  assign _15609_ = \bapg_rd.w_ptr_r [3] ? _15608_ : _15601_;
  assign _15610_ = \bapg_rd.w_ptr_r [4] ? _15609_ : _15594_;
  assign _15611_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [14] : \MSYNC_1r1w.synth.nz.mem[224] [14];
  assign _15612_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [14] : \MSYNC_1r1w.synth.nz.mem[226] [14];
  assign _15613_ = \bapg_rd.w_ptr_r [1] ? _15612_ : _15611_;
  assign _15614_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [14] : \MSYNC_1r1w.synth.nz.mem[228] [14];
  assign _15615_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [14] : \MSYNC_1r1w.synth.nz.mem[230] [14];
  assign _15616_ = \bapg_rd.w_ptr_r [1] ? _15615_ : _15614_;
  assign _15617_ = \bapg_rd.w_ptr_r [2] ? _15616_ : _15613_;
  assign _15618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [14] : \MSYNC_1r1w.synth.nz.mem[232] [14];
  assign _15619_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [14] : \MSYNC_1r1w.synth.nz.mem[234] [14];
  assign _15620_ = \bapg_rd.w_ptr_r [1] ? _15619_ : _15618_;
  assign _15621_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [14] : \MSYNC_1r1w.synth.nz.mem[236] [14];
  assign _15622_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [14] : \MSYNC_1r1w.synth.nz.mem[238] [14];
  assign _15623_ = \bapg_rd.w_ptr_r [1] ? _15622_ : _15621_;
  assign _15624_ = \bapg_rd.w_ptr_r [2] ? _15623_ : _15620_;
  assign _15625_ = \bapg_rd.w_ptr_r [3] ? _15624_ : _15617_;
  assign _15626_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [14] : \MSYNC_1r1w.synth.nz.mem[240] [14];
  assign _15627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [14] : \MSYNC_1r1w.synth.nz.mem[242] [14];
  assign _15628_ = \bapg_rd.w_ptr_r [1] ? _15627_ : _15626_;
  assign _15629_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [14] : \MSYNC_1r1w.synth.nz.mem[244] [14];
  assign _15630_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [14] : \MSYNC_1r1w.synth.nz.mem[246] [14];
  assign _15631_ = \bapg_rd.w_ptr_r [1] ? _15630_ : _15629_;
  assign _15632_ = \bapg_rd.w_ptr_r [2] ? _15631_ : _15628_;
  assign _15633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [14] : \MSYNC_1r1w.synth.nz.mem[248] [14];
  assign _15634_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [14] : \MSYNC_1r1w.synth.nz.mem[250] [14];
  assign _15635_ = \bapg_rd.w_ptr_r [1] ? _15634_ : _15633_;
  assign _15636_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [14] : \MSYNC_1r1w.synth.nz.mem[252] [14];
  assign _15637_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [14] : \MSYNC_1r1w.synth.nz.mem[254] [14];
  assign _15638_ = \bapg_rd.w_ptr_r [1] ? _15637_ : _15636_;
  assign _15639_ = \bapg_rd.w_ptr_r [2] ? _15638_ : _15635_;
  assign _15640_ = \bapg_rd.w_ptr_r [3] ? _15639_ : _15632_;
  assign _15641_ = \bapg_rd.w_ptr_r [4] ? _15640_ : _15625_;
  assign _15642_ = \bapg_rd.w_ptr_r [5] ? _15641_ : _15610_;
  assign _15643_ = \bapg_rd.w_ptr_r [6] ? _15642_ : _15579_;
  assign _15644_ = \bapg_rd.w_ptr_r [7] ? _15643_ : _15516_;
  assign _15645_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [14] : \MSYNC_1r1w.synth.nz.mem[256] [14];
  assign _15646_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [14] : \MSYNC_1r1w.synth.nz.mem[258] [14];
  assign _15647_ = \bapg_rd.w_ptr_r [1] ? _15646_ : _15645_;
  assign _15648_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [14] : \MSYNC_1r1w.synth.nz.mem[260] [14];
  assign _15649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [14] : \MSYNC_1r1w.synth.nz.mem[262] [14];
  assign _15650_ = \bapg_rd.w_ptr_r [1] ? _15649_ : _15648_;
  assign _15651_ = \bapg_rd.w_ptr_r [2] ? _15650_ : _15647_;
  assign _15652_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [14] : \MSYNC_1r1w.synth.nz.mem[264] [14];
  assign _15653_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [14] : \MSYNC_1r1w.synth.nz.mem[266] [14];
  assign _15654_ = \bapg_rd.w_ptr_r [1] ? _15653_ : _15652_;
  assign _15655_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [14] : \MSYNC_1r1w.synth.nz.mem[268] [14];
  assign _15656_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [14] : \MSYNC_1r1w.synth.nz.mem[270] [14];
  assign _15657_ = \bapg_rd.w_ptr_r [1] ? _15656_ : _15655_;
  assign _15658_ = \bapg_rd.w_ptr_r [2] ? _15657_ : _15654_;
  assign _15659_ = \bapg_rd.w_ptr_r [3] ? _15658_ : _15651_;
  assign _15660_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [14] : \MSYNC_1r1w.synth.nz.mem[272] [14];
  assign _15661_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [14] : \MSYNC_1r1w.synth.nz.mem[274] [14];
  assign _15662_ = \bapg_rd.w_ptr_r [1] ? _15661_ : _15660_;
  assign _15663_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [14] : \MSYNC_1r1w.synth.nz.mem[276] [14];
  assign _15664_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [14] : \MSYNC_1r1w.synth.nz.mem[278] [14];
  assign _15665_ = \bapg_rd.w_ptr_r [1] ? _15664_ : _15663_;
  assign _15666_ = \bapg_rd.w_ptr_r [2] ? _15665_ : _15662_;
  assign _15667_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [14] : \MSYNC_1r1w.synth.nz.mem[280] [14];
  assign _15668_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [14] : \MSYNC_1r1w.synth.nz.mem[282] [14];
  assign _15669_ = \bapg_rd.w_ptr_r [1] ? _15668_ : _15667_;
  assign _15670_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [14] : \MSYNC_1r1w.synth.nz.mem[284] [14];
  assign _15671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [14] : \MSYNC_1r1w.synth.nz.mem[286] [14];
  assign _15672_ = \bapg_rd.w_ptr_r [1] ? _15671_ : _15670_;
  assign _15673_ = \bapg_rd.w_ptr_r [2] ? _15672_ : _15669_;
  assign _15674_ = \bapg_rd.w_ptr_r [3] ? _15673_ : _15666_;
  assign _15675_ = \bapg_rd.w_ptr_r [4] ? _15674_ : _15659_;
  assign _15676_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [14] : \MSYNC_1r1w.synth.nz.mem[288] [14];
  assign _15677_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [14] : \MSYNC_1r1w.synth.nz.mem[290] [14];
  assign _15678_ = \bapg_rd.w_ptr_r [1] ? _15677_ : _15676_;
  assign _15679_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [14] : \MSYNC_1r1w.synth.nz.mem[292] [14];
  assign _15680_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [14] : \MSYNC_1r1w.synth.nz.mem[294] [14];
  assign _15681_ = \bapg_rd.w_ptr_r [1] ? _15680_ : _15679_;
  assign _15682_ = \bapg_rd.w_ptr_r [2] ? _15681_ : _15678_;
  assign _15683_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [14] : \MSYNC_1r1w.synth.nz.mem[296] [14];
  assign _15684_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [14] : \MSYNC_1r1w.synth.nz.mem[298] [14];
  assign _15685_ = \bapg_rd.w_ptr_r [1] ? _15684_ : _15683_;
  assign _15686_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [14] : \MSYNC_1r1w.synth.nz.mem[300] [14];
  assign _15687_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [14] : \MSYNC_1r1w.synth.nz.mem[302] [14];
  assign _15688_ = \bapg_rd.w_ptr_r [1] ? _15687_ : _15686_;
  assign _15689_ = \bapg_rd.w_ptr_r [2] ? _15688_ : _15685_;
  assign _15690_ = \bapg_rd.w_ptr_r [3] ? _15689_ : _15682_;
  assign _15691_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [14] : \MSYNC_1r1w.synth.nz.mem[304] [14];
  assign _15692_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [14] : \MSYNC_1r1w.synth.nz.mem[306] [14];
  assign _15693_ = \bapg_rd.w_ptr_r [1] ? _15692_ : _15691_;
  assign _15694_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [14] : \MSYNC_1r1w.synth.nz.mem[308] [14];
  assign _15695_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [14] : \MSYNC_1r1w.synth.nz.mem[310] [14];
  assign _15696_ = \bapg_rd.w_ptr_r [1] ? _15695_ : _15694_;
  assign _15697_ = \bapg_rd.w_ptr_r [2] ? _15696_ : _15693_;
  assign _15698_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [14] : \MSYNC_1r1w.synth.nz.mem[312] [14];
  assign _15699_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [14] : \MSYNC_1r1w.synth.nz.mem[314] [14];
  assign _15700_ = \bapg_rd.w_ptr_r [1] ? _15699_ : _15698_;
  assign _15701_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [14] : \MSYNC_1r1w.synth.nz.mem[316] [14];
  assign _15702_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [14] : \MSYNC_1r1w.synth.nz.mem[318] [14];
  assign _15703_ = \bapg_rd.w_ptr_r [1] ? _15702_ : _15701_;
  assign _15704_ = \bapg_rd.w_ptr_r [2] ? _15703_ : _15700_;
  assign _15705_ = \bapg_rd.w_ptr_r [3] ? _15704_ : _15697_;
  assign _15706_ = \bapg_rd.w_ptr_r [4] ? _15705_ : _15690_;
  assign _15707_ = \bapg_rd.w_ptr_r [5] ? _15706_ : _15675_;
  assign _15708_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [14] : \MSYNC_1r1w.synth.nz.mem[320] [14];
  assign _15709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [14] : \MSYNC_1r1w.synth.nz.mem[322] [14];
  assign _15710_ = \bapg_rd.w_ptr_r [1] ? _15709_ : _15708_;
  assign _15711_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [14] : \MSYNC_1r1w.synth.nz.mem[324] [14];
  assign _15712_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [14] : \MSYNC_1r1w.synth.nz.mem[326] [14];
  assign _15713_ = \bapg_rd.w_ptr_r [1] ? _15712_ : _15711_;
  assign _15714_ = \bapg_rd.w_ptr_r [2] ? _15713_ : _15710_;
  assign _15715_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [14] : \MSYNC_1r1w.synth.nz.mem[328] [14];
  assign _15716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [14] : \MSYNC_1r1w.synth.nz.mem[330] [14];
  assign _15717_ = \bapg_rd.w_ptr_r [1] ? _15716_ : _15715_;
  assign _15718_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [14] : \MSYNC_1r1w.synth.nz.mem[332] [14];
  assign _15719_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [14] : \MSYNC_1r1w.synth.nz.mem[334] [14];
  assign _15720_ = \bapg_rd.w_ptr_r [1] ? _15719_ : _15718_;
  assign _15721_ = \bapg_rd.w_ptr_r [2] ? _15720_ : _15717_;
  assign _15722_ = \bapg_rd.w_ptr_r [3] ? _15721_ : _15714_;
  assign _15723_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [14] : \MSYNC_1r1w.synth.nz.mem[336] [14];
  assign _15724_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [14] : \MSYNC_1r1w.synth.nz.mem[338] [14];
  assign _15725_ = \bapg_rd.w_ptr_r [1] ? _15724_ : _15723_;
  assign _15726_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [14] : \MSYNC_1r1w.synth.nz.mem[340] [14];
  assign _15727_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [14] : \MSYNC_1r1w.synth.nz.mem[342] [14];
  assign _15728_ = \bapg_rd.w_ptr_r [1] ? _15727_ : _15726_;
  assign _15729_ = \bapg_rd.w_ptr_r [2] ? _15728_ : _15725_;
  assign _15730_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [14] : \MSYNC_1r1w.synth.nz.mem[344] [14];
  assign _15731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [14] : \MSYNC_1r1w.synth.nz.mem[346] [14];
  assign _15732_ = \bapg_rd.w_ptr_r [1] ? _15731_ : _15730_;
  assign _15733_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [14] : \MSYNC_1r1w.synth.nz.mem[348] [14];
  assign _15734_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [14] : \MSYNC_1r1w.synth.nz.mem[350] [14];
  assign _15735_ = \bapg_rd.w_ptr_r [1] ? _15734_ : _15733_;
  assign _15736_ = \bapg_rd.w_ptr_r [2] ? _15735_ : _15732_;
  assign _15737_ = \bapg_rd.w_ptr_r [3] ? _15736_ : _15729_;
  assign _15738_ = \bapg_rd.w_ptr_r [4] ? _15737_ : _15722_;
  assign _15739_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [14] : \MSYNC_1r1w.synth.nz.mem[352] [14];
  assign _15740_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [14] : \MSYNC_1r1w.synth.nz.mem[354] [14];
  assign _15741_ = \bapg_rd.w_ptr_r [1] ? _15740_ : _15739_;
  assign _15742_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [14] : \MSYNC_1r1w.synth.nz.mem[356] [14];
  assign _15743_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [14] : \MSYNC_1r1w.synth.nz.mem[358] [14];
  assign _15744_ = \bapg_rd.w_ptr_r [1] ? _15743_ : _15742_;
  assign _15745_ = \bapg_rd.w_ptr_r [2] ? _15744_ : _15741_;
  assign _15746_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [14] : \MSYNC_1r1w.synth.nz.mem[360] [14];
  assign _15747_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [14] : \MSYNC_1r1w.synth.nz.mem[362] [14];
  assign _15748_ = \bapg_rd.w_ptr_r [1] ? _15747_ : _15746_;
  assign _15749_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [14] : \MSYNC_1r1w.synth.nz.mem[364] [14];
  assign _15750_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [14] : \MSYNC_1r1w.synth.nz.mem[366] [14];
  assign _15751_ = \bapg_rd.w_ptr_r [1] ? _15750_ : _15749_;
  assign _15752_ = \bapg_rd.w_ptr_r [2] ? _15751_ : _15748_;
  assign _15753_ = \bapg_rd.w_ptr_r [3] ? _15752_ : _15745_;
  assign _15754_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [14] : \MSYNC_1r1w.synth.nz.mem[368] [14];
  assign _15755_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [14] : \MSYNC_1r1w.synth.nz.mem[370] [14];
  assign _15756_ = \bapg_rd.w_ptr_r [1] ? _15755_ : _15754_;
  assign _15757_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [14] : \MSYNC_1r1w.synth.nz.mem[372] [14];
  assign _15758_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [14] : \MSYNC_1r1w.synth.nz.mem[374] [14];
  assign _15759_ = \bapg_rd.w_ptr_r [1] ? _15758_ : _15757_;
  assign _15760_ = \bapg_rd.w_ptr_r [2] ? _15759_ : _15756_;
  assign _15761_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [14] : \MSYNC_1r1w.synth.nz.mem[376] [14];
  assign _15762_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [14] : \MSYNC_1r1w.synth.nz.mem[378] [14];
  assign _15763_ = \bapg_rd.w_ptr_r [1] ? _15762_ : _15761_;
  assign _15764_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [14] : \MSYNC_1r1w.synth.nz.mem[380] [14];
  assign _15765_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [14] : \MSYNC_1r1w.synth.nz.mem[382] [14];
  assign _15766_ = \bapg_rd.w_ptr_r [1] ? _15765_ : _15764_;
  assign _15767_ = \bapg_rd.w_ptr_r [2] ? _15766_ : _15763_;
  assign _15768_ = \bapg_rd.w_ptr_r [3] ? _15767_ : _15760_;
  assign _15769_ = \bapg_rd.w_ptr_r [4] ? _15768_ : _15753_;
  assign _15770_ = \bapg_rd.w_ptr_r [5] ? _15769_ : _15738_;
  assign _15771_ = \bapg_rd.w_ptr_r [6] ? _15770_ : _15707_;
  assign _15772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [14] : \MSYNC_1r1w.synth.nz.mem[384] [14];
  assign _15773_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [14] : \MSYNC_1r1w.synth.nz.mem[386] [14];
  assign _15774_ = \bapg_rd.w_ptr_r [1] ? _15773_ : _15772_;
  assign _15775_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [14] : \MSYNC_1r1w.synth.nz.mem[388] [14];
  assign _15776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [14] : \MSYNC_1r1w.synth.nz.mem[390] [14];
  assign _15777_ = \bapg_rd.w_ptr_r [1] ? _15776_ : _15775_;
  assign _15778_ = \bapg_rd.w_ptr_r [2] ? _15777_ : _15774_;
  assign _15779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [14] : \MSYNC_1r1w.synth.nz.mem[392] [14];
  assign _15780_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [14] : \MSYNC_1r1w.synth.nz.mem[394] [14];
  assign _15781_ = \bapg_rd.w_ptr_r [1] ? _15780_ : _15779_;
  assign _15782_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [14] : \MSYNC_1r1w.synth.nz.mem[396] [14];
  assign _15783_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [14] : \MSYNC_1r1w.synth.nz.mem[398] [14];
  assign _15784_ = \bapg_rd.w_ptr_r [1] ? _15783_ : _15782_;
  assign _15785_ = \bapg_rd.w_ptr_r [2] ? _15784_ : _15781_;
  assign _15786_ = \bapg_rd.w_ptr_r [3] ? _15785_ : _15778_;
  assign _15787_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [14] : \MSYNC_1r1w.synth.nz.mem[400] [14];
  assign _15788_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [14] : \MSYNC_1r1w.synth.nz.mem[402] [14];
  assign _15789_ = \bapg_rd.w_ptr_r [1] ? _15788_ : _15787_;
  assign _15790_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [14] : \MSYNC_1r1w.synth.nz.mem[404] [14];
  assign _15791_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [14] : \MSYNC_1r1w.synth.nz.mem[406] [14];
  assign _15792_ = \bapg_rd.w_ptr_r [1] ? _15791_ : _15790_;
  assign _15793_ = \bapg_rd.w_ptr_r [2] ? _15792_ : _15789_;
  assign _15794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [14] : \MSYNC_1r1w.synth.nz.mem[408] [14];
  assign _15795_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [14] : \MSYNC_1r1w.synth.nz.mem[410] [14];
  assign _15796_ = \bapg_rd.w_ptr_r [1] ? _15795_ : _15794_;
  assign _15797_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [14] : \MSYNC_1r1w.synth.nz.mem[412] [14];
  assign _15798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [14] : \MSYNC_1r1w.synth.nz.mem[414] [14];
  assign _15799_ = \bapg_rd.w_ptr_r [1] ? _15798_ : _15797_;
  assign _15800_ = \bapg_rd.w_ptr_r [2] ? _15799_ : _15796_;
  assign _15801_ = \bapg_rd.w_ptr_r [3] ? _15800_ : _15793_;
  assign _15802_ = \bapg_rd.w_ptr_r [4] ? _15801_ : _15786_;
  assign _15803_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [14] : \MSYNC_1r1w.synth.nz.mem[416] [14];
  assign _15804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [14] : \MSYNC_1r1w.synth.nz.mem[418] [14];
  assign _15805_ = \bapg_rd.w_ptr_r [1] ? _15804_ : _15803_;
  assign _15806_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [14] : \MSYNC_1r1w.synth.nz.mem[420] [14];
  assign _15807_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [14] : \MSYNC_1r1w.synth.nz.mem[422] [14];
  assign _15808_ = \bapg_rd.w_ptr_r [1] ? _15807_ : _15806_;
  assign _15809_ = \bapg_rd.w_ptr_r [2] ? _15808_ : _15805_;
  assign _15810_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [14] : \MSYNC_1r1w.synth.nz.mem[424] [14];
  assign _15811_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [14] : \MSYNC_1r1w.synth.nz.mem[426] [14];
  assign _15812_ = \bapg_rd.w_ptr_r [1] ? _15811_ : _15810_;
  assign _15813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [14] : \MSYNC_1r1w.synth.nz.mem[428] [14];
  assign _15814_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [14] : \MSYNC_1r1w.synth.nz.mem[430] [14];
  assign _15815_ = \bapg_rd.w_ptr_r [1] ? _15814_ : _15813_;
  assign _15816_ = \bapg_rd.w_ptr_r [2] ? _15815_ : _15812_;
  assign _15817_ = \bapg_rd.w_ptr_r [3] ? _15816_ : _15809_;
  assign _15818_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [14] : \MSYNC_1r1w.synth.nz.mem[432] [14];
  assign _15819_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [14] : \MSYNC_1r1w.synth.nz.mem[434] [14];
  assign _15820_ = \bapg_rd.w_ptr_r [1] ? _15819_ : _15818_;
  assign _15821_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [14] : \MSYNC_1r1w.synth.nz.mem[436] [14];
  assign _15822_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [14] : \MSYNC_1r1w.synth.nz.mem[438] [14];
  assign _15823_ = \bapg_rd.w_ptr_r [1] ? _15822_ : _15821_;
  assign _15824_ = \bapg_rd.w_ptr_r [2] ? _15823_ : _15820_;
  assign _15825_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [14] : \MSYNC_1r1w.synth.nz.mem[440] [14];
  assign _15826_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [14] : \MSYNC_1r1w.synth.nz.mem[442] [14];
  assign _15827_ = \bapg_rd.w_ptr_r [1] ? _15826_ : _15825_;
  assign _15828_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [14] : \MSYNC_1r1w.synth.nz.mem[444] [14];
  assign _15829_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [14] : \MSYNC_1r1w.synth.nz.mem[446] [14];
  assign _15830_ = \bapg_rd.w_ptr_r [1] ? _15829_ : _15828_;
  assign _15831_ = \bapg_rd.w_ptr_r [2] ? _15830_ : _15827_;
  assign _15832_ = \bapg_rd.w_ptr_r [3] ? _15831_ : _15824_;
  assign _15833_ = \bapg_rd.w_ptr_r [4] ? _15832_ : _15817_;
  assign _15834_ = \bapg_rd.w_ptr_r [5] ? _15833_ : _15802_;
  assign _15835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [14] : \MSYNC_1r1w.synth.nz.mem[448] [14];
  assign _15836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [14] : \MSYNC_1r1w.synth.nz.mem[450] [14];
  assign _15837_ = \bapg_rd.w_ptr_r [1] ? _15836_ : _15835_;
  assign _15838_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [14] : \MSYNC_1r1w.synth.nz.mem[452] [14];
  assign _15839_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [14] : \MSYNC_1r1w.synth.nz.mem[454] [14];
  assign _15840_ = \bapg_rd.w_ptr_r [1] ? _15839_ : _15838_;
  assign _15841_ = \bapg_rd.w_ptr_r [2] ? _15840_ : _15837_;
  assign _15842_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [14] : \MSYNC_1r1w.synth.nz.mem[456] [14];
  assign _15843_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [14] : \MSYNC_1r1w.synth.nz.mem[458] [14];
  assign _15844_ = \bapg_rd.w_ptr_r [1] ? _15843_ : _15842_;
  assign _15845_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [14] : \MSYNC_1r1w.synth.nz.mem[460] [14];
  assign _15846_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [14] : \MSYNC_1r1w.synth.nz.mem[462] [14];
  assign _15847_ = \bapg_rd.w_ptr_r [1] ? _15846_ : _15845_;
  assign _15848_ = \bapg_rd.w_ptr_r [2] ? _15847_ : _15844_;
  assign _15849_ = \bapg_rd.w_ptr_r [3] ? _15848_ : _15841_;
  assign _15850_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [14] : \MSYNC_1r1w.synth.nz.mem[464] [14];
  assign _15851_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [14] : \MSYNC_1r1w.synth.nz.mem[466] [14];
  assign _15852_ = \bapg_rd.w_ptr_r [1] ? _15851_ : _15850_;
  assign _15853_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [14] : \MSYNC_1r1w.synth.nz.mem[468] [14];
  assign _15854_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [14] : \MSYNC_1r1w.synth.nz.mem[470] [14];
  assign _15855_ = \bapg_rd.w_ptr_r [1] ? _15854_ : _15853_;
  assign _15856_ = \bapg_rd.w_ptr_r [2] ? _15855_ : _15852_;
  assign _15857_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [14] : \MSYNC_1r1w.synth.nz.mem[472] [14];
  assign _15858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [14] : \MSYNC_1r1w.synth.nz.mem[474] [14];
  assign _15859_ = \bapg_rd.w_ptr_r [1] ? _15858_ : _15857_;
  assign _15860_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [14] : \MSYNC_1r1w.synth.nz.mem[476] [14];
  assign _15861_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [14] : \MSYNC_1r1w.synth.nz.mem[478] [14];
  assign _15862_ = \bapg_rd.w_ptr_r [1] ? _15861_ : _15860_;
  assign _15863_ = \bapg_rd.w_ptr_r [2] ? _15862_ : _15859_;
  assign _15864_ = \bapg_rd.w_ptr_r [3] ? _15863_ : _15856_;
  assign _15865_ = \bapg_rd.w_ptr_r [4] ? _15864_ : _15849_;
  assign _15866_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [14] : \MSYNC_1r1w.synth.nz.mem[480] [14];
  assign _15867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [14] : \MSYNC_1r1w.synth.nz.mem[482] [14];
  assign _15868_ = \bapg_rd.w_ptr_r [1] ? _15867_ : _15866_;
  assign _15869_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [14] : \MSYNC_1r1w.synth.nz.mem[484] [14];
  assign _15870_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [14] : \MSYNC_1r1w.synth.nz.mem[486] [14];
  assign _15871_ = \bapg_rd.w_ptr_r [1] ? _15870_ : _15869_;
  assign _15872_ = \bapg_rd.w_ptr_r [2] ? _15871_ : _15868_;
  assign _15873_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [14] : \MSYNC_1r1w.synth.nz.mem[488] [14];
  assign _15874_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [14] : \MSYNC_1r1w.synth.nz.mem[490] [14];
  assign _15875_ = \bapg_rd.w_ptr_r [1] ? _15874_ : _15873_;
  assign _15876_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [14] : \MSYNC_1r1w.synth.nz.mem[492] [14];
  assign _15877_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [14] : \MSYNC_1r1w.synth.nz.mem[494] [14];
  assign _15878_ = \bapg_rd.w_ptr_r [1] ? _15877_ : _15876_;
  assign _15879_ = \bapg_rd.w_ptr_r [2] ? _15878_ : _15875_;
  assign _15880_ = \bapg_rd.w_ptr_r [3] ? _15879_ : _15872_;
  assign _15881_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [14] : \MSYNC_1r1w.synth.nz.mem[496] [14];
  assign _15882_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [14] : \MSYNC_1r1w.synth.nz.mem[498] [14];
  assign _15883_ = \bapg_rd.w_ptr_r [1] ? _15882_ : _15881_;
  assign _15884_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [14] : \MSYNC_1r1w.synth.nz.mem[500] [14];
  assign _15885_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [14] : \MSYNC_1r1w.synth.nz.mem[502] [14];
  assign _15886_ = \bapg_rd.w_ptr_r [1] ? _15885_ : _15884_;
  assign _15887_ = \bapg_rd.w_ptr_r [2] ? _15886_ : _15883_;
  assign _15888_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [14] : \MSYNC_1r1w.synth.nz.mem[504] [14];
  assign _15889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [14] : \MSYNC_1r1w.synth.nz.mem[506] [14];
  assign _15890_ = \bapg_rd.w_ptr_r [1] ? _15889_ : _15888_;
  assign _15891_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [14] : \MSYNC_1r1w.synth.nz.mem[508] [14];
  assign _15892_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [14] : \MSYNC_1r1w.synth.nz.mem[510] [14];
  assign _15893_ = \bapg_rd.w_ptr_r [1] ? _15892_ : _15891_;
  assign _15894_ = \bapg_rd.w_ptr_r [2] ? _15893_ : _15890_;
  assign _15895_ = \bapg_rd.w_ptr_r [3] ? _15894_ : _15887_;
  assign _15896_ = \bapg_rd.w_ptr_r [4] ? _15895_ : _15880_;
  assign _15897_ = \bapg_rd.w_ptr_r [5] ? _15896_ : _15865_;
  assign _15898_ = \bapg_rd.w_ptr_r [6] ? _15897_ : _15834_;
  assign _15899_ = \bapg_rd.w_ptr_r [7] ? _15898_ : _15771_;
  assign _15900_ = \bapg_rd.w_ptr_r [8] ? _15899_ : _15644_;
  assign _15901_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [14] : \MSYNC_1r1w.synth.nz.mem[512] [14];
  assign _15902_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [14] : \MSYNC_1r1w.synth.nz.mem[514] [14];
  assign _15903_ = \bapg_rd.w_ptr_r [1] ? _15902_ : _15901_;
  assign _15904_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [14] : \MSYNC_1r1w.synth.nz.mem[516] [14];
  assign _15905_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [14] : \MSYNC_1r1w.synth.nz.mem[518] [14];
  assign _15906_ = \bapg_rd.w_ptr_r [1] ? _15905_ : _15904_;
  assign _15907_ = \bapg_rd.w_ptr_r [2] ? _15906_ : _15903_;
  assign _15908_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [14] : \MSYNC_1r1w.synth.nz.mem[520] [14];
  assign _15909_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [14] : \MSYNC_1r1w.synth.nz.mem[522] [14];
  assign _15910_ = \bapg_rd.w_ptr_r [1] ? _15909_ : _15908_;
  assign _15911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [14] : \MSYNC_1r1w.synth.nz.mem[524] [14];
  assign _15912_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [14] : \MSYNC_1r1w.synth.nz.mem[526] [14];
  assign _15913_ = \bapg_rd.w_ptr_r [1] ? _15912_ : _15911_;
  assign _15914_ = \bapg_rd.w_ptr_r [2] ? _15913_ : _15910_;
  assign _15915_ = \bapg_rd.w_ptr_r [3] ? _15914_ : _15907_;
  assign _15916_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [14] : \MSYNC_1r1w.synth.nz.mem[528] [14];
  assign _15917_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [14] : \MSYNC_1r1w.synth.nz.mem[530] [14];
  assign _15918_ = \bapg_rd.w_ptr_r [1] ? _15917_ : _15916_;
  assign _15919_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [14] : \MSYNC_1r1w.synth.nz.mem[532] [14];
  assign _15920_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [14] : \MSYNC_1r1w.synth.nz.mem[534] [14];
  assign _15921_ = \bapg_rd.w_ptr_r [1] ? _15920_ : _15919_;
  assign _15922_ = \bapg_rd.w_ptr_r [2] ? _15921_ : _15918_;
  assign _15923_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [14] : \MSYNC_1r1w.synth.nz.mem[536] [14];
  assign _15924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [14] : \MSYNC_1r1w.synth.nz.mem[538] [14];
  assign _15925_ = \bapg_rd.w_ptr_r [1] ? _15924_ : _15923_;
  assign _15926_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [14] : \MSYNC_1r1w.synth.nz.mem[540] [14];
  assign _15927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [14] : \MSYNC_1r1w.synth.nz.mem[542] [14];
  assign _15928_ = \bapg_rd.w_ptr_r [1] ? _15927_ : _15926_;
  assign _15929_ = \bapg_rd.w_ptr_r [2] ? _15928_ : _15925_;
  assign _15930_ = \bapg_rd.w_ptr_r [3] ? _15929_ : _15922_;
  assign _15931_ = \bapg_rd.w_ptr_r [4] ? _15930_ : _15915_;
  assign _15932_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [14] : \MSYNC_1r1w.synth.nz.mem[544] [14];
  assign _15933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [14] : \MSYNC_1r1w.synth.nz.mem[546] [14];
  assign _15934_ = \bapg_rd.w_ptr_r [1] ? _15933_ : _15932_;
  assign _15935_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [14] : \MSYNC_1r1w.synth.nz.mem[548] [14];
  assign _15936_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [14] : \MSYNC_1r1w.synth.nz.mem[550] [14];
  assign _15937_ = \bapg_rd.w_ptr_r [1] ? _15936_ : _15935_;
  assign _15938_ = \bapg_rd.w_ptr_r [2] ? _15937_ : _15934_;
  assign _15939_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [14] : \MSYNC_1r1w.synth.nz.mem[552] [14];
  assign _15940_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [14] : \MSYNC_1r1w.synth.nz.mem[554] [14];
  assign _15941_ = \bapg_rd.w_ptr_r [1] ? _15940_ : _15939_;
  assign _15942_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [14] : \MSYNC_1r1w.synth.nz.mem[556] [14];
  assign _15943_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [14] : \MSYNC_1r1w.synth.nz.mem[558] [14];
  assign _15944_ = \bapg_rd.w_ptr_r [1] ? _15943_ : _15942_;
  assign _15945_ = \bapg_rd.w_ptr_r [2] ? _15944_ : _15941_;
  assign _15946_ = \bapg_rd.w_ptr_r [3] ? _15945_ : _15938_;
  assign _15947_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [14] : \MSYNC_1r1w.synth.nz.mem[560] [14];
  assign _15948_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [14] : \MSYNC_1r1w.synth.nz.mem[562] [14];
  assign _15949_ = \bapg_rd.w_ptr_r [1] ? _15948_ : _15947_;
  assign _15950_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [14] : \MSYNC_1r1w.synth.nz.mem[564] [14];
  assign _15951_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [14] : \MSYNC_1r1w.synth.nz.mem[566] [14];
  assign _15952_ = \bapg_rd.w_ptr_r [1] ? _15951_ : _15950_;
  assign _15953_ = \bapg_rd.w_ptr_r [2] ? _15952_ : _15949_;
  assign _15954_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [14] : \MSYNC_1r1w.synth.nz.mem[568] [14];
  assign _15955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [14] : \MSYNC_1r1w.synth.nz.mem[570] [14];
  assign _15956_ = \bapg_rd.w_ptr_r [1] ? _15955_ : _15954_;
  assign _15957_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [14] : \MSYNC_1r1w.synth.nz.mem[572] [14];
  assign _15958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [14] : \MSYNC_1r1w.synth.nz.mem[574] [14];
  assign _15959_ = \bapg_rd.w_ptr_r [1] ? _15958_ : _15957_;
  assign _15960_ = \bapg_rd.w_ptr_r [2] ? _15959_ : _15956_;
  assign _15961_ = \bapg_rd.w_ptr_r [3] ? _15960_ : _15953_;
  assign _15962_ = \bapg_rd.w_ptr_r [4] ? _15961_ : _15946_;
  assign _15963_ = \bapg_rd.w_ptr_r [5] ? _15962_ : _15931_;
  assign _15964_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [14] : \MSYNC_1r1w.synth.nz.mem[576] [14];
  assign _15965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [14] : \MSYNC_1r1w.synth.nz.mem[578] [14];
  assign _15966_ = \bapg_rd.w_ptr_r [1] ? _15965_ : _15964_;
  assign _15967_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [14] : \MSYNC_1r1w.synth.nz.mem[580] [14];
  assign _15968_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [14] : \MSYNC_1r1w.synth.nz.mem[582] [14];
  assign _15969_ = \bapg_rd.w_ptr_r [1] ? _15968_ : _15967_;
  assign _15970_ = \bapg_rd.w_ptr_r [2] ? _15969_ : _15966_;
  assign _15971_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [14] : \MSYNC_1r1w.synth.nz.mem[584] [14];
  assign _15972_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [14] : \MSYNC_1r1w.synth.nz.mem[586] [14];
  assign _15973_ = \bapg_rd.w_ptr_r [1] ? _15972_ : _15971_;
  assign _15974_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [14] : \MSYNC_1r1w.synth.nz.mem[588] [14];
  assign _15975_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [14] : \MSYNC_1r1w.synth.nz.mem[590] [14];
  assign _15976_ = \bapg_rd.w_ptr_r [1] ? _15975_ : _15974_;
  assign _15977_ = \bapg_rd.w_ptr_r [2] ? _15976_ : _15973_;
  assign _15978_ = \bapg_rd.w_ptr_r [3] ? _15977_ : _15970_;
  assign _15979_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [14] : \MSYNC_1r1w.synth.nz.mem[592] [14];
  assign _15980_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [14] : \MSYNC_1r1w.synth.nz.mem[594] [14];
  assign _15981_ = \bapg_rd.w_ptr_r [1] ? _15980_ : _15979_;
  assign _15982_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [14] : \MSYNC_1r1w.synth.nz.mem[596] [14];
  assign _15983_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [14] : \MSYNC_1r1w.synth.nz.mem[598] [14];
  assign _15984_ = \bapg_rd.w_ptr_r [1] ? _15983_ : _15982_;
  assign _15985_ = \bapg_rd.w_ptr_r [2] ? _15984_ : _15981_;
  assign _15986_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [14] : \MSYNC_1r1w.synth.nz.mem[600] [14];
  assign _15987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [14] : \MSYNC_1r1w.synth.nz.mem[602] [14];
  assign _15988_ = \bapg_rd.w_ptr_r [1] ? _15987_ : _15986_;
  assign _15989_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [14] : \MSYNC_1r1w.synth.nz.mem[604] [14];
  assign _15990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [14] : \MSYNC_1r1w.synth.nz.mem[606] [14];
  assign _15991_ = \bapg_rd.w_ptr_r [1] ? _15990_ : _15989_;
  assign _15992_ = \bapg_rd.w_ptr_r [2] ? _15991_ : _15988_;
  assign _15993_ = \bapg_rd.w_ptr_r [3] ? _15992_ : _15985_;
  assign _15994_ = \bapg_rd.w_ptr_r [4] ? _15993_ : _15978_;
  assign _15995_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [14] : \MSYNC_1r1w.synth.nz.mem[608] [14];
  assign _15996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [14] : \MSYNC_1r1w.synth.nz.mem[610] [14];
  assign _15997_ = \bapg_rd.w_ptr_r [1] ? _15996_ : _15995_;
  assign _15998_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [14] : \MSYNC_1r1w.synth.nz.mem[612] [14];
  assign _15999_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [14] : \MSYNC_1r1w.synth.nz.mem[614] [14];
  assign _16000_ = \bapg_rd.w_ptr_r [1] ? _15999_ : _15998_;
  assign _16001_ = \bapg_rd.w_ptr_r [2] ? _16000_ : _15997_;
  assign _16002_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [14] : \MSYNC_1r1w.synth.nz.mem[616] [14];
  assign _16003_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [14] : \MSYNC_1r1w.synth.nz.mem[618] [14];
  assign _16004_ = \bapg_rd.w_ptr_r [1] ? _16003_ : _16002_;
  assign _16005_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [14] : \MSYNC_1r1w.synth.nz.mem[620] [14];
  assign _16006_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [14] : \MSYNC_1r1w.synth.nz.mem[622] [14];
  assign _16007_ = \bapg_rd.w_ptr_r [1] ? _16006_ : _16005_;
  assign _16008_ = \bapg_rd.w_ptr_r [2] ? _16007_ : _16004_;
  assign _16009_ = \bapg_rd.w_ptr_r [3] ? _16008_ : _16001_;
  assign _16010_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [14] : \MSYNC_1r1w.synth.nz.mem[624] [14];
  assign _16011_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [14] : \MSYNC_1r1w.synth.nz.mem[626] [14];
  assign _16012_ = \bapg_rd.w_ptr_r [1] ? _16011_ : _16010_;
  assign _16013_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [14] : \MSYNC_1r1w.synth.nz.mem[628] [14];
  assign _16014_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [14] : \MSYNC_1r1w.synth.nz.mem[630] [14];
  assign _16015_ = \bapg_rd.w_ptr_r [1] ? _16014_ : _16013_;
  assign _16016_ = \bapg_rd.w_ptr_r [2] ? _16015_ : _16012_;
  assign _16017_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [14] : \MSYNC_1r1w.synth.nz.mem[632] [14];
  assign _16018_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [14] : \MSYNC_1r1w.synth.nz.mem[634] [14];
  assign _16019_ = \bapg_rd.w_ptr_r [1] ? _16018_ : _16017_;
  assign _16020_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [14] : \MSYNC_1r1w.synth.nz.mem[636] [14];
  assign _16021_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [14] : \MSYNC_1r1w.synth.nz.mem[638] [14];
  assign _16022_ = \bapg_rd.w_ptr_r [1] ? _16021_ : _16020_;
  assign _16023_ = \bapg_rd.w_ptr_r [2] ? _16022_ : _16019_;
  assign _16024_ = \bapg_rd.w_ptr_r [3] ? _16023_ : _16016_;
  assign _16025_ = \bapg_rd.w_ptr_r [4] ? _16024_ : _16009_;
  assign _16026_ = \bapg_rd.w_ptr_r [5] ? _16025_ : _15994_;
  assign _16027_ = \bapg_rd.w_ptr_r [6] ? _16026_ : _15963_;
  assign _16028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [14] : \MSYNC_1r1w.synth.nz.mem[640] [14];
  assign _16029_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [14] : \MSYNC_1r1w.synth.nz.mem[642] [14];
  assign _16030_ = \bapg_rd.w_ptr_r [1] ? _16029_ : _16028_;
  assign _16031_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [14] : \MSYNC_1r1w.synth.nz.mem[644] [14];
  assign _16032_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [14] : \MSYNC_1r1w.synth.nz.mem[646] [14];
  assign _16033_ = \bapg_rd.w_ptr_r [1] ? _16032_ : _16031_;
  assign _16034_ = \bapg_rd.w_ptr_r [2] ? _16033_ : _16030_;
  assign _16035_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [14] : \MSYNC_1r1w.synth.nz.mem[648] [14];
  assign _16036_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [14] : \MSYNC_1r1w.synth.nz.mem[650] [14];
  assign _16037_ = \bapg_rd.w_ptr_r [1] ? _16036_ : _16035_;
  assign _16038_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [14] : \MSYNC_1r1w.synth.nz.mem[652] [14];
  assign _16039_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [14] : \MSYNC_1r1w.synth.nz.mem[654] [14];
  assign _16040_ = \bapg_rd.w_ptr_r [1] ? _16039_ : _16038_;
  assign _16041_ = \bapg_rd.w_ptr_r [2] ? _16040_ : _16037_;
  assign _16042_ = \bapg_rd.w_ptr_r [3] ? _16041_ : _16034_;
  assign _16043_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [14] : \MSYNC_1r1w.synth.nz.mem[656] [14];
  assign _16044_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [14] : \MSYNC_1r1w.synth.nz.mem[658] [14];
  assign _16045_ = \bapg_rd.w_ptr_r [1] ? _16044_ : _16043_;
  assign _16046_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [14] : \MSYNC_1r1w.synth.nz.mem[660] [14];
  assign _16047_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [14] : \MSYNC_1r1w.synth.nz.mem[662] [14];
  assign _16048_ = \bapg_rd.w_ptr_r [1] ? _16047_ : _16046_;
  assign _16049_ = \bapg_rd.w_ptr_r [2] ? _16048_ : _16045_;
  assign _16050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [14] : \MSYNC_1r1w.synth.nz.mem[664] [14];
  assign _16051_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [14] : \MSYNC_1r1w.synth.nz.mem[666] [14];
  assign _16052_ = \bapg_rd.w_ptr_r [1] ? _16051_ : _16050_;
  assign _16053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [14] : \MSYNC_1r1w.synth.nz.mem[668] [14];
  assign _16054_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [14] : \MSYNC_1r1w.synth.nz.mem[670] [14];
  assign _16055_ = \bapg_rd.w_ptr_r [1] ? _16054_ : _16053_;
  assign _16056_ = \bapg_rd.w_ptr_r [2] ? _16055_ : _16052_;
  assign _16057_ = \bapg_rd.w_ptr_r [3] ? _16056_ : _16049_;
  assign _16058_ = \bapg_rd.w_ptr_r [4] ? _16057_ : _16042_;
  assign _16059_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [14] : \MSYNC_1r1w.synth.nz.mem[672] [14];
  assign _16060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [14] : \MSYNC_1r1w.synth.nz.mem[674] [14];
  assign _16061_ = \bapg_rd.w_ptr_r [1] ? _16060_ : _16059_;
  assign _16062_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [14] : \MSYNC_1r1w.synth.nz.mem[676] [14];
  assign _16063_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [14] : \MSYNC_1r1w.synth.nz.mem[678] [14];
  assign _16064_ = \bapg_rd.w_ptr_r [1] ? _16063_ : _16062_;
  assign _16065_ = \bapg_rd.w_ptr_r [2] ? _16064_ : _16061_;
  assign _16066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [14] : \MSYNC_1r1w.synth.nz.mem[680] [14];
  assign _16067_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [14] : \MSYNC_1r1w.synth.nz.mem[682] [14];
  assign _16068_ = \bapg_rd.w_ptr_r [1] ? _16067_ : _16066_;
  assign _16069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [14] : \MSYNC_1r1w.synth.nz.mem[684] [14];
  assign _16070_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [14] : \MSYNC_1r1w.synth.nz.mem[686] [14];
  assign _16071_ = \bapg_rd.w_ptr_r [1] ? _16070_ : _16069_;
  assign _16072_ = \bapg_rd.w_ptr_r [2] ? _16071_ : _16068_;
  assign _16073_ = \bapg_rd.w_ptr_r [3] ? _16072_ : _16065_;
  assign _16074_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [14] : \MSYNC_1r1w.synth.nz.mem[688] [14];
  assign _16075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [14] : \MSYNC_1r1w.synth.nz.mem[690] [14];
  assign _16076_ = \bapg_rd.w_ptr_r [1] ? _16075_ : _16074_;
  assign _16077_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [14] : \MSYNC_1r1w.synth.nz.mem[692] [14];
  assign _16078_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [14] : \MSYNC_1r1w.synth.nz.mem[694] [14];
  assign _16079_ = \bapg_rd.w_ptr_r [1] ? _16078_ : _16077_;
  assign _16080_ = \bapg_rd.w_ptr_r [2] ? _16079_ : _16076_;
  assign _16081_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [14] : \MSYNC_1r1w.synth.nz.mem[696] [14];
  assign _16082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [14] : \MSYNC_1r1w.synth.nz.mem[698] [14];
  assign _16083_ = \bapg_rd.w_ptr_r [1] ? _16082_ : _16081_;
  assign _16084_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [14] : \MSYNC_1r1w.synth.nz.mem[700] [14];
  assign _16085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [14] : \MSYNC_1r1w.synth.nz.mem[702] [14];
  assign _16086_ = \bapg_rd.w_ptr_r [1] ? _16085_ : _16084_;
  assign _16087_ = \bapg_rd.w_ptr_r [2] ? _16086_ : _16083_;
  assign _16088_ = \bapg_rd.w_ptr_r [3] ? _16087_ : _16080_;
  assign _16089_ = \bapg_rd.w_ptr_r [4] ? _16088_ : _16073_;
  assign _16090_ = \bapg_rd.w_ptr_r [5] ? _16089_ : _16058_;
  assign _16091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [14] : \MSYNC_1r1w.synth.nz.mem[704] [14];
  assign _16092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [14] : \MSYNC_1r1w.synth.nz.mem[706] [14];
  assign _16093_ = \bapg_rd.w_ptr_r [1] ? _16092_ : _16091_;
  assign _16094_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [14] : \MSYNC_1r1w.synth.nz.mem[708] [14];
  assign _16095_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [14] : \MSYNC_1r1w.synth.nz.mem[710] [14];
  assign _16096_ = \bapg_rd.w_ptr_r [1] ? _16095_ : _16094_;
  assign _16097_ = \bapg_rd.w_ptr_r [2] ? _16096_ : _16093_;
  assign _16098_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [14] : \MSYNC_1r1w.synth.nz.mem[712] [14];
  assign _16099_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [14] : \MSYNC_1r1w.synth.nz.mem[714] [14];
  assign _16100_ = \bapg_rd.w_ptr_r [1] ? _16099_ : _16098_;
  assign _16101_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [14] : \MSYNC_1r1w.synth.nz.mem[716] [14];
  assign _16102_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [14] : \MSYNC_1r1w.synth.nz.mem[718] [14];
  assign _16103_ = \bapg_rd.w_ptr_r [1] ? _16102_ : _16101_;
  assign _16104_ = \bapg_rd.w_ptr_r [2] ? _16103_ : _16100_;
  assign _16105_ = \bapg_rd.w_ptr_r [3] ? _16104_ : _16097_;
  assign _16106_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [14] : \MSYNC_1r1w.synth.nz.mem[720] [14];
  assign _16107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [14] : \MSYNC_1r1w.synth.nz.mem[722] [14];
  assign _16108_ = \bapg_rd.w_ptr_r [1] ? _16107_ : _16106_;
  assign _16109_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [14] : \MSYNC_1r1w.synth.nz.mem[724] [14];
  assign _16110_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [14] : \MSYNC_1r1w.synth.nz.mem[726] [14];
  assign _16111_ = \bapg_rd.w_ptr_r [1] ? _16110_ : _16109_;
  assign _16112_ = \bapg_rd.w_ptr_r [2] ? _16111_ : _16108_;
  assign _16113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [14] : \MSYNC_1r1w.synth.nz.mem[728] [14];
  assign _16114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [14] : \MSYNC_1r1w.synth.nz.mem[730] [14];
  assign _16115_ = \bapg_rd.w_ptr_r [1] ? _16114_ : _16113_;
  assign _16116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [14] : \MSYNC_1r1w.synth.nz.mem[732] [14];
  assign _16117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [14] : \MSYNC_1r1w.synth.nz.mem[734] [14];
  assign _16118_ = \bapg_rd.w_ptr_r [1] ? _16117_ : _16116_;
  assign _16119_ = \bapg_rd.w_ptr_r [2] ? _16118_ : _16115_;
  assign _16120_ = \bapg_rd.w_ptr_r [3] ? _16119_ : _16112_;
  assign _16121_ = \bapg_rd.w_ptr_r [4] ? _16120_ : _16105_;
  assign _16122_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [14] : \MSYNC_1r1w.synth.nz.mem[736] [14];
  assign _16123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [14] : \MSYNC_1r1w.synth.nz.mem[738] [14];
  assign _16124_ = \bapg_rd.w_ptr_r [1] ? _16123_ : _16122_;
  assign _16125_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [14] : \MSYNC_1r1w.synth.nz.mem[740] [14];
  assign _16126_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [14] : \MSYNC_1r1w.synth.nz.mem[742] [14];
  assign _16127_ = \bapg_rd.w_ptr_r [1] ? _16126_ : _16125_;
  assign _16128_ = \bapg_rd.w_ptr_r [2] ? _16127_ : _16124_;
  assign _16129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [14] : \MSYNC_1r1w.synth.nz.mem[744] [14];
  assign _16130_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [14] : \MSYNC_1r1w.synth.nz.mem[746] [14];
  assign _16131_ = \bapg_rd.w_ptr_r [1] ? _16130_ : _16129_;
  assign _16132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [14] : \MSYNC_1r1w.synth.nz.mem[748] [14];
  assign _16133_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [14] : \MSYNC_1r1w.synth.nz.mem[750] [14];
  assign _16134_ = \bapg_rd.w_ptr_r [1] ? _16133_ : _16132_;
  assign _16135_ = \bapg_rd.w_ptr_r [2] ? _16134_ : _16131_;
  assign _16136_ = \bapg_rd.w_ptr_r [3] ? _16135_ : _16128_;
  assign _16137_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [14] : \MSYNC_1r1w.synth.nz.mem[752] [14];
  assign _16138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [14] : \MSYNC_1r1w.synth.nz.mem[754] [14];
  assign _16139_ = \bapg_rd.w_ptr_r [1] ? _16138_ : _16137_;
  assign _16140_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [14] : \MSYNC_1r1w.synth.nz.mem[756] [14];
  assign _16141_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [14] : \MSYNC_1r1w.synth.nz.mem[758] [14];
  assign _16142_ = \bapg_rd.w_ptr_r [1] ? _16141_ : _16140_;
  assign _16143_ = \bapg_rd.w_ptr_r [2] ? _16142_ : _16139_;
  assign _16144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [14] : \MSYNC_1r1w.synth.nz.mem[760] [14];
  assign _16145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [14] : \MSYNC_1r1w.synth.nz.mem[762] [14];
  assign _16146_ = \bapg_rd.w_ptr_r [1] ? _16145_ : _16144_;
  assign _16147_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [14] : \MSYNC_1r1w.synth.nz.mem[764] [14];
  assign _16148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [14] : \MSYNC_1r1w.synth.nz.mem[766] [14];
  assign _16149_ = \bapg_rd.w_ptr_r [1] ? _16148_ : _16147_;
  assign _16150_ = \bapg_rd.w_ptr_r [2] ? _16149_ : _16146_;
  assign _16151_ = \bapg_rd.w_ptr_r [3] ? _16150_ : _16143_;
  assign _16152_ = \bapg_rd.w_ptr_r [4] ? _16151_ : _16136_;
  assign _16153_ = \bapg_rd.w_ptr_r [5] ? _16152_ : _16121_;
  assign _16154_ = \bapg_rd.w_ptr_r [6] ? _16153_ : _16090_;
  assign _16155_ = \bapg_rd.w_ptr_r [7] ? _16154_ : _16027_;
  assign _16156_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [14] : \MSYNC_1r1w.synth.nz.mem[768] [14];
  assign _16157_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [14] : \MSYNC_1r1w.synth.nz.mem[770] [14];
  assign _16158_ = \bapg_rd.w_ptr_r [1] ? _16157_ : _16156_;
  assign _16159_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [14] : \MSYNC_1r1w.synth.nz.mem[772] [14];
  assign _16160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [14] : \MSYNC_1r1w.synth.nz.mem[774] [14];
  assign _16161_ = \bapg_rd.w_ptr_r [1] ? _16160_ : _16159_;
  assign _16162_ = \bapg_rd.w_ptr_r [2] ? _16161_ : _16158_;
  assign _16163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [14] : \MSYNC_1r1w.synth.nz.mem[776] [14];
  assign _16164_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [14] : \MSYNC_1r1w.synth.nz.mem[778] [14];
  assign _16165_ = \bapg_rd.w_ptr_r [1] ? _16164_ : _16163_;
  assign _16166_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [14] : \MSYNC_1r1w.synth.nz.mem[780] [14];
  assign _16167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [14] : \MSYNC_1r1w.synth.nz.mem[782] [14];
  assign _16168_ = \bapg_rd.w_ptr_r [1] ? _16167_ : _16166_;
  assign _16169_ = \bapg_rd.w_ptr_r [2] ? _16168_ : _16165_;
  assign _16170_ = \bapg_rd.w_ptr_r [3] ? _16169_ : _16162_;
  assign _16171_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [14] : \MSYNC_1r1w.synth.nz.mem[784] [14];
  assign _16172_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [14] : \MSYNC_1r1w.synth.nz.mem[786] [14];
  assign _16173_ = \bapg_rd.w_ptr_r [1] ? _16172_ : _16171_;
  assign _16174_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [14] : \MSYNC_1r1w.synth.nz.mem[788] [14];
  assign _16175_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [14] : \MSYNC_1r1w.synth.nz.mem[790] [14];
  assign _16176_ = \bapg_rd.w_ptr_r [1] ? _16175_ : _16174_;
  assign _16177_ = \bapg_rd.w_ptr_r [2] ? _16176_ : _16173_;
  assign _16178_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [14] : \MSYNC_1r1w.synth.nz.mem[792] [14];
  assign _16179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [14] : \MSYNC_1r1w.synth.nz.mem[794] [14];
  assign _16180_ = \bapg_rd.w_ptr_r [1] ? _16179_ : _16178_;
  assign _16181_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [14] : \MSYNC_1r1w.synth.nz.mem[796] [14];
  assign _16182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [14] : \MSYNC_1r1w.synth.nz.mem[798] [14];
  assign _16183_ = \bapg_rd.w_ptr_r [1] ? _16182_ : _16181_;
  assign _16184_ = \bapg_rd.w_ptr_r [2] ? _16183_ : _16180_;
  assign _16185_ = \bapg_rd.w_ptr_r [3] ? _16184_ : _16177_;
  assign _16186_ = \bapg_rd.w_ptr_r [4] ? _16185_ : _16170_;
  assign _16187_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [14] : \MSYNC_1r1w.synth.nz.mem[800] [14];
  assign _16188_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [14] : \MSYNC_1r1w.synth.nz.mem[802] [14];
  assign _16189_ = \bapg_rd.w_ptr_r [1] ? _16188_ : _16187_;
  assign _16190_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [14] : \MSYNC_1r1w.synth.nz.mem[804] [14];
  assign _16191_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [14] : \MSYNC_1r1w.synth.nz.mem[806] [14];
  assign _16192_ = \bapg_rd.w_ptr_r [1] ? _16191_ : _16190_;
  assign _16193_ = \bapg_rd.w_ptr_r [2] ? _16192_ : _16189_;
  assign _16194_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [14] : \MSYNC_1r1w.synth.nz.mem[808] [14];
  assign _16195_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [14] : \MSYNC_1r1w.synth.nz.mem[810] [14];
  assign _16196_ = \bapg_rd.w_ptr_r [1] ? _16195_ : _16194_;
  assign _16197_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [14] : \MSYNC_1r1w.synth.nz.mem[812] [14];
  assign _16198_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [14] : \MSYNC_1r1w.synth.nz.mem[814] [14];
  assign _16199_ = \bapg_rd.w_ptr_r [1] ? _16198_ : _16197_;
  assign _16200_ = \bapg_rd.w_ptr_r [2] ? _16199_ : _16196_;
  assign _16201_ = \bapg_rd.w_ptr_r [3] ? _16200_ : _16193_;
  assign _16202_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [14] : \MSYNC_1r1w.synth.nz.mem[816] [14];
  assign _16203_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [14] : \MSYNC_1r1w.synth.nz.mem[818] [14];
  assign _16204_ = \bapg_rd.w_ptr_r [1] ? _16203_ : _16202_;
  assign _16205_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [14] : \MSYNC_1r1w.synth.nz.mem[820] [14];
  assign _16206_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [14] : \MSYNC_1r1w.synth.nz.mem[822] [14];
  assign _16207_ = \bapg_rd.w_ptr_r [1] ? _16206_ : _16205_;
  assign _16208_ = \bapg_rd.w_ptr_r [2] ? _16207_ : _16204_;
  assign _16209_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [14] : \MSYNC_1r1w.synth.nz.mem[824] [14];
  assign _16210_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [14] : \MSYNC_1r1w.synth.nz.mem[826] [14];
  assign _16211_ = \bapg_rd.w_ptr_r [1] ? _16210_ : _16209_;
  assign _16212_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [14] : \MSYNC_1r1w.synth.nz.mem[828] [14];
  assign _16213_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [14] : \MSYNC_1r1w.synth.nz.mem[830] [14];
  assign _16214_ = \bapg_rd.w_ptr_r [1] ? _16213_ : _16212_;
  assign _16215_ = \bapg_rd.w_ptr_r [2] ? _16214_ : _16211_;
  assign _16216_ = \bapg_rd.w_ptr_r [3] ? _16215_ : _16208_;
  assign _16217_ = \bapg_rd.w_ptr_r [4] ? _16216_ : _16201_;
  assign _16218_ = \bapg_rd.w_ptr_r [5] ? _16217_ : _16186_;
  assign _16219_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [14] : \MSYNC_1r1w.synth.nz.mem[832] [14];
  assign _16220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [14] : \MSYNC_1r1w.synth.nz.mem[834] [14];
  assign _16221_ = \bapg_rd.w_ptr_r [1] ? _16220_ : _16219_;
  assign _16222_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [14] : \MSYNC_1r1w.synth.nz.mem[836] [14];
  assign _16223_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [14] : \MSYNC_1r1w.synth.nz.mem[838] [14];
  assign _16224_ = \bapg_rd.w_ptr_r [1] ? _16223_ : _16222_;
  assign _16225_ = \bapg_rd.w_ptr_r [2] ? _16224_ : _16221_;
  assign _16226_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [14] : \MSYNC_1r1w.synth.nz.mem[840] [14];
  assign _16227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [14] : \MSYNC_1r1w.synth.nz.mem[842] [14];
  assign _16228_ = \bapg_rd.w_ptr_r [1] ? _16227_ : _16226_;
  assign _16229_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [14] : \MSYNC_1r1w.synth.nz.mem[844] [14];
  assign _16230_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [14] : \MSYNC_1r1w.synth.nz.mem[846] [14];
  assign _16231_ = \bapg_rd.w_ptr_r [1] ? _16230_ : _16229_;
  assign _16232_ = \bapg_rd.w_ptr_r [2] ? _16231_ : _16228_;
  assign _16233_ = \bapg_rd.w_ptr_r [3] ? _16232_ : _16225_;
  assign _16234_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [14] : \MSYNC_1r1w.synth.nz.mem[848] [14];
  assign _16235_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [14] : \MSYNC_1r1w.synth.nz.mem[850] [14];
  assign _16236_ = \bapg_rd.w_ptr_r [1] ? _16235_ : _16234_;
  assign _16237_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [14] : \MSYNC_1r1w.synth.nz.mem[852] [14];
  assign _16238_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [14] : \MSYNC_1r1w.synth.nz.mem[854] [14];
  assign _16239_ = \bapg_rd.w_ptr_r [1] ? _16238_ : _16237_;
  assign _16240_ = \bapg_rd.w_ptr_r [2] ? _16239_ : _16236_;
  assign _16241_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [14] : \MSYNC_1r1w.synth.nz.mem[856] [14];
  assign _16242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [14] : \MSYNC_1r1w.synth.nz.mem[858] [14];
  assign _16243_ = \bapg_rd.w_ptr_r [1] ? _16242_ : _16241_;
  assign _16244_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [14] : \MSYNC_1r1w.synth.nz.mem[860] [14];
  assign _16245_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [14] : \MSYNC_1r1w.synth.nz.mem[862] [14];
  assign _16246_ = \bapg_rd.w_ptr_r [1] ? _16245_ : _16244_;
  assign _16247_ = \bapg_rd.w_ptr_r [2] ? _16246_ : _16243_;
  assign _16248_ = \bapg_rd.w_ptr_r [3] ? _16247_ : _16240_;
  assign _16249_ = \bapg_rd.w_ptr_r [4] ? _16248_ : _16233_;
  assign _16250_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [14] : \MSYNC_1r1w.synth.nz.mem[864] [14];
  assign _16251_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [14] : \MSYNC_1r1w.synth.nz.mem[866] [14];
  assign _16252_ = \bapg_rd.w_ptr_r [1] ? _16251_ : _16250_;
  assign _16253_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [14] : \MSYNC_1r1w.synth.nz.mem[868] [14];
  assign _16254_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [14] : \MSYNC_1r1w.synth.nz.mem[870] [14];
  assign _16255_ = \bapg_rd.w_ptr_r [1] ? _16254_ : _16253_;
  assign _16256_ = \bapg_rd.w_ptr_r [2] ? _16255_ : _16252_;
  assign _16257_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [14] : \MSYNC_1r1w.synth.nz.mem[872] [14];
  assign _16258_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [14] : \MSYNC_1r1w.synth.nz.mem[874] [14];
  assign _16259_ = \bapg_rd.w_ptr_r [1] ? _16258_ : _16257_;
  assign _16260_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [14] : \MSYNC_1r1w.synth.nz.mem[876] [14];
  assign _16261_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [14] : \MSYNC_1r1w.synth.nz.mem[878] [14];
  assign _16262_ = \bapg_rd.w_ptr_r [1] ? _16261_ : _16260_;
  assign _16263_ = \bapg_rd.w_ptr_r [2] ? _16262_ : _16259_;
  assign _16264_ = \bapg_rd.w_ptr_r [3] ? _16263_ : _16256_;
  assign _16265_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [14] : \MSYNC_1r1w.synth.nz.mem[880] [14];
  assign _16266_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [14] : \MSYNC_1r1w.synth.nz.mem[882] [14];
  assign _16267_ = \bapg_rd.w_ptr_r [1] ? _16266_ : _16265_;
  assign _16268_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [14] : \MSYNC_1r1w.synth.nz.mem[884] [14];
  assign _16269_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [14] : \MSYNC_1r1w.synth.nz.mem[886] [14];
  assign _16270_ = \bapg_rd.w_ptr_r [1] ? _16269_ : _16268_;
  assign _16271_ = \bapg_rd.w_ptr_r [2] ? _16270_ : _16267_;
  assign _16272_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [14] : \MSYNC_1r1w.synth.nz.mem[888] [14];
  assign _16273_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [14] : \MSYNC_1r1w.synth.nz.mem[890] [14];
  assign _16274_ = \bapg_rd.w_ptr_r [1] ? _16273_ : _16272_;
  assign _16275_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [14] : \MSYNC_1r1w.synth.nz.mem[892] [14];
  assign _16276_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [14] : \MSYNC_1r1w.synth.nz.mem[894] [14];
  assign _16277_ = \bapg_rd.w_ptr_r [1] ? _16276_ : _16275_;
  assign _16278_ = \bapg_rd.w_ptr_r [2] ? _16277_ : _16274_;
  assign _16279_ = \bapg_rd.w_ptr_r [3] ? _16278_ : _16271_;
  assign _16280_ = \bapg_rd.w_ptr_r [4] ? _16279_ : _16264_;
  assign _16281_ = \bapg_rd.w_ptr_r [5] ? _16280_ : _16249_;
  assign _16282_ = \bapg_rd.w_ptr_r [6] ? _16281_ : _16218_;
  assign _16283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [14] : \MSYNC_1r1w.synth.nz.mem[896] [14];
  assign _16284_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [14] : \MSYNC_1r1w.synth.nz.mem[898] [14];
  assign _16285_ = \bapg_rd.w_ptr_r [1] ? _16284_ : _16283_;
  assign _16286_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [14] : \MSYNC_1r1w.synth.nz.mem[900] [14];
  assign _16287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [14] : \MSYNC_1r1w.synth.nz.mem[902] [14];
  assign _16288_ = \bapg_rd.w_ptr_r [1] ? _16287_ : _16286_;
  assign _16289_ = \bapg_rd.w_ptr_r [2] ? _16288_ : _16285_;
  assign _16290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [14] : \MSYNC_1r1w.synth.nz.mem[904] [14];
  assign _16291_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [14] : \MSYNC_1r1w.synth.nz.mem[906] [14];
  assign _16292_ = \bapg_rd.w_ptr_r [1] ? _16291_ : _16290_;
  assign _16293_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [14] : \MSYNC_1r1w.synth.nz.mem[908] [14];
  assign _16294_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [14] : \MSYNC_1r1w.synth.nz.mem[910] [14];
  assign _16295_ = \bapg_rd.w_ptr_r [1] ? _16294_ : _16293_;
  assign _16296_ = \bapg_rd.w_ptr_r [2] ? _16295_ : _16292_;
  assign _16297_ = \bapg_rd.w_ptr_r [3] ? _16296_ : _16289_;
  assign _16298_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [14] : \MSYNC_1r1w.synth.nz.mem[912] [14];
  assign _16299_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [14] : \MSYNC_1r1w.synth.nz.mem[914] [14];
  assign _16300_ = \bapg_rd.w_ptr_r [1] ? _16299_ : _16298_;
  assign _16301_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [14] : \MSYNC_1r1w.synth.nz.mem[916] [14];
  assign _16302_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [14] : \MSYNC_1r1w.synth.nz.mem[918] [14];
  assign _16303_ = \bapg_rd.w_ptr_r [1] ? _16302_ : _16301_;
  assign _16304_ = \bapg_rd.w_ptr_r [2] ? _16303_ : _16300_;
  assign _16305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [14] : \MSYNC_1r1w.synth.nz.mem[920] [14];
  assign _16306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [14] : \MSYNC_1r1w.synth.nz.mem[922] [14];
  assign _16307_ = \bapg_rd.w_ptr_r [1] ? _16306_ : _16305_;
  assign _16308_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [14] : \MSYNC_1r1w.synth.nz.mem[924] [14];
  assign _16309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [14] : \MSYNC_1r1w.synth.nz.mem[926] [14];
  assign _16310_ = \bapg_rd.w_ptr_r [1] ? _16309_ : _16308_;
  assign _16311_ = \bapg_rd.w_ptr_r [2] ? _16310_ : _16307_;
  assign _16312_ = \bapg_rd.w_ptr_r [3] ? _16311_ : _16304_;
  assign _16313_ = \bapg_rd.w_ptr_r [4] ? _16312_ : _16297_;
  assign _16314_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [14] : \MSYNC_1r1w.synth.nz.mem[928] [14];
  assign _16315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [14] : \MSYNC_1r1w.synth.nz.mem[930] [14];
  assign _16316_ = \bapg_rd.w_ptr_r [1] ? _16315_ : _16314_;
  assign _16317_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [14] : \MSYNC_1r1w.synth.nz.mem[932] [14];
  assign _16318_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [14] : \MSYNC_1r1w.synth.nz.mem[934] [14];
  assign _16319_ = \bapg_rd.w_ptr_r [1] ? _16318_ : _16317_;
  assign _16320_ = \bapg_rd.w_ptr_r [2] ? _16319_ : _16316_;
  assign _16321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [14] : \MSYNC_1r1w.synth.nz.mem[936] [14];
  assign _16322_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [14] : \MSYNC_1r1w.synth.nz.mem[938] [14];
  assign _16323_ = \bapg_rd.w_ptr_r [1] ? _16322_ : _16321_;
  assign _16324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [14] : \MSYNC_1r1w.synth.nz.mem[940] [14];
  assign _16325_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [14] : \MSYNC_1r1w.synth.nz.mem[942] [14];
  assign _16326_ = \bapg_rd.w_ptr_r [1] ? _16325_ : _16324_;
  assign _16327_ = \bapg_rd.w_ptr_r [2] ? _16326_ : _16323_;
  assign _16328_ = \bapg_rd.w_ptr_r [3] ? _16327_ : _16320_;
  assign _16329_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [14] : \MSYNC_1r1w.synth.nz.mem[944] [14];
  assign _16330_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [14] : \MSYNC_1r1w.synth.nz.mem[946] [14];
  assign _16331_ = \bapg_rd.w_ptr_r [1] ? _16330_ : _16329_;
  assign _16332_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [14] : \MSYNC_1r1w.synth.nz.mem[948] [14];
  assign _16333_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [14] : \MSYNC_1r1w.synth.nz.mem[950] [14];
  assign _16334_ = \bapg_rd.w_ptr_r [1] ? _16333_ : _16332_;
  assign _16335_ = \bapg_rd.w_ptr_r [2] ? _16334_ : _16331_;
  assign _16336_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [14] : \MSYNC_1r1w.synth.nz.mem[952] [14];
  assign _16337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [14] : \MSYNC_1r1w.synth.nz.mem[954] [14];
  assign _16338_ = \bapg_rd.w_ptr_r [1] ? _16337_ : _16336_;
  assign _16339_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [14] : \MSYNC_1r1w.synth.nz.mem[956] [14];
  assign _16340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [14] : \MSYNC_1r1w.synth.nz.mem[958] [14];
  assign _16341_ = \bapg_rd.w_ptr_r [1] ? _16340_ : _16339_;
  assign _16342_ = \bapg_rd.w_ptr_r [2] ? _16341_ : _16338_;
  assign _16343_ = \bapg_rd.w_ptr_r [3] ? _16342_ : _16335_;
  assign _16344_ = \bapg_rd.w_ptr_r [4] ? _16343_ : _16328_;
  assign _16345_ = \bapg_rd.w_ptr_r [5] ? _16344_ : _16313_;
  assign _16346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [14] : \MSYNC_1r1w.synth.nz.mem[960] [14];
  assign _16347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [14] : \MSYNC_1r1w.synth.nz.mem[962] [14];
  assign _16348_ = \bapg_rd.w_ptr_r [1] ? _16347_ : _16346_;
  assign _16349_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [14] : \MSYNC_1r1w.synth.nz.mem[964] [14];
  assign _16350_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [14] : \MSYNC_1r1w.synth.nz.mem[966] [14];
  assign _16351_ = \bapg_rd.w_ptr_r [1] ? _16350_ : _16349_;
  assign _16352_ = \bapg_rd.w_ptr_r [2] ? _16351_ : _16348_;
  assign _16353_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [14] : \MSYNC_1r1w.synth.nz.mem[968] [14];
  assign _16354_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [14] : \MSYNC_1r1w.synth.nz.mem[970] [14];
  assign _16355_ = \bapg_rd.w_ptr_r [1] ? _16354_ : _16353_;
  assign _16356_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [14] : \MSYNC_1r1w.synth.nz.mem[972] [14];
  assign _16357_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [14] : \MSYNC_1r1w.synth.nz.mem[974] [14];
  assign _16358_ = \bapg_rd.w_ptr_r [1] ? _16357_ : _16356_;
  assign _16359_ = \bapg_rd.w_ptr_r [2] ? _16358_ : _16355_;
  assign _16360_ = \bapg_rd.w_ptr_r [3] ? _16359_ : _16352_;
  assign _16361_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [14] : \MSYNC_1r1w.synth.nz.mem[976] [14];
  assign _16362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [14] : \MSYNC_1r1w.synth.nz.mem[978] [14];
  assign _16363_ = \bapg_rd.w_ptr_r [1] ? _16362_ : _16361_;
  assign _16364_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [14] : \MSYNC_1r1w.synth.nz.mem[980] [14];
  assign _16365_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [14] : \MSYNC_1r1w.synth.nz.mem[982] [14];
  assign _16366_ = \bapg_rd.w_ptr_r [1] ? _16365_ : _16364_;
  assign _16367_ = \bapg_rd.w_ptr_r [2] ? _16366_ : _16363_;
  assign _16368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [14] : \MSYNC_1r1w.synth.nz.mem[984] [14];
  assign _16369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [14] : \MSYNC_1r1w.synth.nz.mem[986] [14];
  assign _16370_ = \bapg_rd.w_ptr_r [1] ? _16369_ : _16368_;
  assign _16371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [14] : \MSYNC_1r1w.synth.nz.mem[988] [14];
  assign _16372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [14] : \MSYNC_1r1w.synth.nz.mem[990] [14];
  assign _16373_ = \bapg_rd.w_ptr_r [1] ? _16372_ : _16371_;
  assign _16374_ = \bapg_rd.w_ptr_r [2] ? _16373_ : _16370_;
  assign _16375_ = \bapg_rd.w_ptr_r [3] ? _16374_ : _16367_;
  assign _16376_ = \bapg_rd.w_ptr_r [4] ? _16375_ : _16360_;
  assign _16377_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [14] : \MSYNC_1r1w.synth.nz.mem[992] [14];
  assign _16378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [14] : \MSYNC_1r1w.synth.nz.mem[994] [14];
  assign _16379_ = \bapg_rd.w_ptr_r [1] ? _16378_ : _16377_;
  assign _16380_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [14] : \MSYNC_1r1w.synth.nz.mem[996] [14];
  assign _16381_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [14] : \MSYNC_1r1w.synth.nz.mem[998] [14];
  assign _16382_ = \bapg_rd.w_ptr_r [1] ? _16381_ : _16380_;
  assign _16383_ = \bapg_rd.w_ptr_r [2] ? _16382_ : _16379_;
  assign _16384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [14] : \MSYNC_1r1w.synth.nz.mem[1000] [14];
  assign _16385_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [14] : \MSYNC_1r1w.synth.nz.mem[1002] [14];
  assign _16386_ = \bapg_rd.w_ptr_r [1] ? _16385_ : _16384_;
  assign _16387_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [14] : \MSYNC_1r1w.synth.nz.mem[1004] [14];
  assign _16388_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [14] : \MSYNC_1r1w.synth.nz.mem[1006] [14];
  assign _16389_ = \bapg_rd.w_ptr_r [1] ? _16388_ : _16387_;
  assign _16390_ = \bapg_rd.w_ptr_r [2] ? _16389_ : _16386_;
  assign _16391_ = \bapg_rd.w_ptr_r [3] ? _16390_ : _16383_;
  assign _16392_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [14] : \MSYNC_1r1w.synth.nz.mem[1008] [14];
  assign _16393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [14] : \MSYNC_1r1w.synth.nz.mem[1010] [14];
  assign _16394_ = \bapg_rd.w_ptr_r [1] ? _16393_ : _16392_;
  assign _16395_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [14] : \MSYNC_1r1w.synth.nz.mem[1012] [14];
  assign _16396_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [14] : \MSYNC_1r1w.synth.nz.mem[1014] [14];
  assign _16397_ = \bapg_rd.w_ptr_r [1] ? _16396_ : _16395_;
  assign _16398_ = \bapg_rd.w_ptr_r [2] ? _16397_ : _16394_;
  assign _16399_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [14] : \MSYNC_1r1w.synth.nz.mem[1016] [14];
  assign _16400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [14] : \MSYNC_1r1w.synth.nz.mem[1018] [14];
  assign _16401_ = \bapg_rd.w_ptr_r [1] ? _16400_ : _16399_;
  assign _16402_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [14] : \MSYNC_1r1w.synth.nz.mem[1020] [14];
  assign _16403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [14] : \MSYNC_1r1w.synth.nz.mem[1022] [14];
  assign _16404_ = \bapg_rd.w_ptr_r [1] ? _16403_ : _16402_;
  assign _16405_ = \bapg_rd.w_ptr_r [2] ? _16404_ : _16401_;
  assign _16406_ = \bapg_rd.w_ptr_r [3] ? _16405_ : _16398_;
  assign _16407_ = \bapg_rd.w_ptr_r [4] ? _16406_ : _16391_;
  assign _16408_ = \bapg_rd.w_ptr_r [5] ? _16407_ : _16376_;
  assign _16409_ = \bapg_rd.w_ptr_r [6] ? _16408_ : _16345_;
  assign _16410_ = \bapg_rd.w_ptr_r [7] ? _16409_ : _16282_;
  assign _16411_ = \bapg_rd.w_ptr_r [8] ? _16410_ : _16155_;
  assign r_data_o[14] = \bapg_rd.w_ptr_r [9] ? _16411_ : _15900_;
  assign _16412_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1] [15] : \MSYNC_1r1w.synth.nz.mem[0] [15];
  assign _16413_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[3] [15] : \MSYNC_1r1w.synth.nz.mem[2] [15];
  assign _16414_ = \bapg_rd.w_ptr_r [1] ? _16413_ : _16412_;
  assign _16415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[5] [15] : \MSYNC_1r1w.synth.nz.mem[4] [15];
  assign _16416_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[7] [15] : \MSYNC_1r1w.synth.nz.mem[6] [15];
  assign _16417_ = \bapg_rd.w_ptr_r [1] ? _16416_ : _16415_;
  assign _16418_ = \bapg_rd.w_ptr_r [2] ? _16417_ : _16414_;
  assign _16419_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[9] [15] : \MSYNC_1r1w.synth.nz.mem[8] [15];
  assign _16420_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[11] [15] : \MSYNC_1r1w.synth.nz.mem[10] [15];
  assign _16421_ = \bapg_rd.w_ptr_r [1] ? _16420_ : _16419_;
  assign _16422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[13] [15] : \MSYNC_1r1w.synth.nz.mem[12] [15];
  assign _16423_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[15] [15] : \MSYNC_1r1w.synth.nz.mem[14] [15];
  assign _16424_ = \bapg_rd.w_ptr_r [1] ? _16423_ : _16422_;
  assign _16425_ = \bapg_rd.w_ptr_r [2] ? _16424_ : _16421_;
  assign _16426_ = \bapg_rd.w_ptr_r [3] ? _16425_ : _16418_;
  assign _16427_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[17] [15] : \MSYNC_1r1w.synth.nz.mem[16] [15];
  assign _16428_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[19] [15] : \MSYNC_1r1w.synth.nz.mem[18] [15];
  assign _16429_ = \bapg_rd.w_ptr_r [1] ? _16428_ : _16427_;
  assign _16430_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[21] [15] : \MSYNC_1r1w.synth.nz.mem[20] [15];
  assign _16431_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[23] [15] : \MSYNC_1r1w.synth.nz.mem[22] [15];
  assign _16432_ = \bapg_rd.w_ptr_r [1] ? _16431_ : _16430_;
  assign _16433_ = \bapg_rd.w_ptr_r [2] ? _16432_ : _16429_;
  assign _16434_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[25] [15] : \MSYNC_1r1w.synth.nz.mem[24] [15];
  assign _16435_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[27] [15] : \MSYNC_1r1w.synth.nz.mem[26] [15];
  assign _16436_ = \bapg_rd.w_ptr_r [1] ? _16435_ : _16434_;
  assign _16437_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[29] [15] : \MSYNC_1r1w.synth.nz.mem[28] [15];
  assign _16438_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[31] [15] : \MSYNC_1r1w.synth.nz.mem[30] [15];
  assign _16439_ = \bapg_rd.w_ptr_r [1] ? _16438_ : _16437_;
  assign _16440_ = \bapg_rd.w_ptr_r [2] ? _16439_ : _16436_;
  assign _16441_ = \bapg_rd.w_ptr_r [3] ? _16440_ : _16433_;
  assign _16442_ = \bapg_rd.w_ptr_r [4] ? _16441_ : _16426_;
  assign _16443_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[33] [15] : \MSYNC_1r1w.synth.nz.mem[32] [15];
  assign _16444_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[35] [15] : \MSYNC_1r1w.synth.nz.mem[34] [15];
  assign _16445_ = \bapg_rd.w_ptr_r [1] ? _16444_ : _16443_;
  assign _16446_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[37] [15] : \MSYNC_1r1w.synth.nz.mem[36] [15];
  assign _16447_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[39] [15] : \MSYNC_1r1w.synth.nz.mem[38] [15];
  assign _16448_ = \bapg_rd.w_ptr_r [1] ? _16447_ : _16446_;
  assign _16449_ = \bapg_rd.w_ptr_r [2] ? _16448_ : _16445_;
  assign _16450_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[41] [15] : \MSYNC_1r1w.synth.nz.mem[40] [15];
  assign _16451_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[43] [15] : \MSYNC_1r1w.synth.nz.mem[42] [15];
  assign _16452_ = \bapg_rd.w_ptr_r [1] ? _16451_ : _16450_;
  assign _16453_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[45] [15] : \MSYNC_1r1w.synth.nz.mem[44] [15];
  assign _16454_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[47] [15] : \MSYNC_1r1w.synth.nz.mem[46] [15];
  assign _16455_ = \bapg_rd.w_ptr_r [1] ? _16454_ : _16453_;
  assign _16456_ = \bapg_rd.w_ptr_r [2] ? _16455_ : _16452_;
  assign _16457_ = \bapg_rd.w_ptr_r [3] ? _16456_ : _16449_;
  assign _16458_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[49] [15] : \MSYNC_1r1w.synth.nz.mem[48] [15];
  assign _16459_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[51] [15] : \MSYNC_1r1w.synth.nz.mem[50] [15];
  assign _16460_ = \bapg_rd.w_ptr_r [1] ? _16459_ : _16458_;
  assign _16461_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[53] [15] : \MSYNC_1r1w.synth.nz.mem[52] [15];
  assign _16462_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[55] [15] : \MSYNC_1r1w.synth.nz.mem[54] [15];
  assign _16463_ = \bapg_rd.w_ptr_r [1] ? _16462_ : _16461_;
  assign _16464_ = \bapg_rd.w_ptr_r [2] ? _16463_ : _16460_;
  assign _16465_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[57] [15] : \MSYNC_1r1w.synth.nz.mem[56] [15];
  assign _16466_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[59] [15] : \MSYNC_1r1w.synth.nz.mem[58] [15];
  assign _16467_ = \bapg_rd.w_ptr_r [1] ? _16466_ : _16465_;
  assign _16468_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[61] [15] : \MSYNC_1r1w.synth.nz.mem[60] [15];
  assign _16469_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[63] [15] : \MSYNC_1r1w.synth.nz.mem[62] [15];
  assign _16470_ = \bapg_rd.w_ptr_r [1] ? _16469_ : _16468_;
  assign _16471_ = \bapg_rd.w_ptr_r [2] ? _16470_ : _16467_;
  assign _16472_ = \bapg_rd.w_ptr_r [3] ? _16471_ : _16464_;
  assign _16473_ = \bapg_rd.w_ptr_r [4] ? _16472_ : _16457_;
  assign _16474_ = \bapg_rd.w_ptr_r [5] ? _16473_ : _16442_;
  assign _16475_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[65] [15] : \MSYNC_1r1w.synth.nz.mem[64] [15];
  assign _16476_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[67] [15] : \MSYNC_1r1w.synth.nz.mem[66] [15];
  assign _16477_ = \bapg_rd.w_ptr_r [1] ? _16476_ : _16475_;
  assign _16478_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[69] [15] : \MSYNC_1r1w.synth.nz.mem[68] [15];
  assign _16479_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[71] [15] : \MSYNC_1r1w.synth.nz.mem[70] [15];
  assign _16480_ = \bapg_rd.w_ptr_r [1] ? _16479_ : _16478_;
  assign _16481_ = \bapg_rd.w_ptr_r [2] ? _16480_ : _16477_;
  assign _16482_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[73] [15] : \MSYNC_1r1w.synth.nz.mem[72] [15];
  assign _16483_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[75] [15] : \MSYNC_1r1w.synth.nz.mem[74] [15];
  assign _16484_ = \bapg_rd.w_ptr_r [1] ? _16483_ : _16482_;
  assign _16485_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[77] [15] : \MSYNC_1r1w.synth.nz.mem[76] [15];
  assign _16486_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[79] [15] : \MSYNC_1r1w.synth.nz.mem[78] [15];
  assign _16487_ = \bapg_rd.w_ptr_r [1] ? _16486_ : _16485_;
  assign _16488_ = \bapg_rd.w_ptr_r [2] ? _16487_ : _16484_;
  assign _16489_ = \bapg_rd.w_ptr_r [3] ? _16488_ : _16481_;
  assign _16490_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[81] [15] : \MSYNC_1r1w.synth.nz.mem[80] [15];
  assign _16491_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[83] [15] : \MSYNC_1r1w.synth.nz.mem[82] [15];
  assign _16492_ = \bapg_rd.w_ptr_r [1] ? _16491_ : _16490_;
  assign _16493_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[85] [15] : \MSYNC_1r1w.synth.nz.mem[84] [15];
  assign _16494_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[87] [15] : \MSYNC_1r1w.synth.nz.mem[86] [15];
  assign _16495_ = \bapg_rd.w_ptr_r [1] ? _16494_ : _16493_;
  assign _16496_ = \bapg_rd.w_ptr_r [2] ? _16495_ : _16492_;
  assign _16497_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[89] [15] : \MSYNC_1r1w.synth.nz.mem[88] [15];
  assign _16498_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[91] [15] : \MSYNC_1r1w.synth.nz.mem[90] [15];
  assign _16499_ = \bapg_rd.w_ptr_r [1] ? _16498_ : _16497_;
  assign _16500_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[93] [15] : \MSYNC_1r1w.synth.nz.mem[92] [15];
  assign _16501_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[95] [15] : \MSYNC_1r1w.synth.nz.mem[94] [15];
  assign _16502_ = \bapg_rd.w_ptr_r [1] ? _16501_ : _16500_;
  assign _16503_ = \bapg_rd.w_ptr_r [2] ? _16502_ : _16499_;
  assign _16504_ = \bapg_rd.w_ptr_r [3] ? _16503_ : _16496_;
  assign _16505_ = \bapg_rd.w_ptr_r [4] ? _16504_ : _16489_;
  assign _16506_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[97] [15] : \MSYNC_1r1w.synth.nz.mem[96] [15];
  assign _16507_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[99] [15] : \MSYNC_1r1w.synth.nz.mem[98] [15];
  assign _16508_ = \bapg_rd.w_ptr_r [1] ? _16507_ : _16506_;
  assign _16509_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[101] [15] : \MSYNC_1r1w.synth.nz.mem[100] [15];
  assign _16510_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[103] [15] : \MSYNC_1r1w.synth.nz.mem[102] [15];
  assign _16511_ = \bapg_rd.w_ptr_r [1] ? _16510_ : _16509_;
  assign _16512_ = \bapg_rd.w_ptr_r [2] ? _16511_ : _16508_;
  assign _16513_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[105] [15] : \MSYNC_1r1w.synth.nz.mem[104] [15];
  assign _16514_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[107] [15] : \MSYNC_1r1w.synth.nz.mem[106] [15];
  assign _16515_ = \bapg_rd.w_ptr_r [1] ? _16514_ : _16513_;
  assign _16516_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[109] [15] : \MSYNC_1r1w.synth.nz.mem[108] [15];
  assign _16517_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[111] [15] : \MSYNC_1r1w.synth.nz.mem[110] [15];
  assign _16518_ = \bapg_rd.w_ptr_r [1] ? _16517_ : _16516_;
  assign _16519_ = \bapg_rd.w_ptr_r [2] ? _16518_ : _16515_;
  assign _16520_ = \bapg_rd.w_ptr_r [3] ? _16519_ : _16512_;
  assign _16521_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[113] [15] : \MSYNC_1r1w.synth.nz.mem[112] [15];
  assign _16522_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[115] [15] : \MSYNC_1r1w.synth.nz.mem[114] [15];
  assign _16523_ = \bapg_rd.w_ptr_r [1] ? _16522_ : _16521_;
  assign _16524_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[117] [15] : \MSYNC_1r1w.synth.nz.mem[116] [15];
  assign _16525_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[119] [15] : \MSYNC_1r1w.synth.nz.mem[118] [15];
  assign _16526_ = \bapg_rd.w_ptr_r [1] ? _16525_ : _16524_;
  assign _16527_ = \bapg_rd.w_ptr_r [2] ? _16526_ : _16523_;
  assign _16528_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[121] [15] : \MSYNC_1r1w.synth.nz.mem[120] [15];
  assign _16529_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[123] [15] : \MSYNC_1r1w.synth.nz.mem[122] [15];
  assign _16530_ = \bapg_rd.w_ptr_r [1] ? _16529_ : _16528_;
  assign _16531_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[125] [15] : \MSYNC_1r1w.synth.nz.mem[124] [15];
  assign _16532_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[127] [15] : \MSYNC_1r1w.synth.nz.mem[126] [15];
  assign _16533_ = \bapg_rd.w_ptr_r [1] ? _16532_ : _16531_;
  assign _16534_ = \bapg_rd.w_ptr_r [2] ? _16533_ : _16530_;
  assign _16535_ = \bapg_rd.w_ptr_r [3] ? _16534_ : _16527_;
  assign _16536_ = \bapg_rd.w_ptr_r [4] ? _16535_ : _16520_;
  assign _16537_ = \bapg_rd.w_ptr_r [5] ? _16536_ : _16505_;
  assign _16538_ = \bapg_rd.w_ptr_r [6] ? _16537_ : _16474_;
  assign _16539_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[129] [15] : \MSYNC_1r1w.synth.nz.mem[128] [15];
  assign _16540_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[131] [15] : \MSYNC_1r1w.synth.nz.mem[130] [15];
  assign _16541_ = \bapg_rd.w_ptr_r [1] ? _16540_ : _16539_;
  assign _16542_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[133] [15] : \MSYNC_1r1w.synth.nz.mem[132] [15];
  assign _16543_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[135] [15] : \MSYNC_1r1w.synth.nz.mem[134] [15];
  assign _16544_ = \bapg_rd.w_ptr_r [1] ? _16543_ : _16542_;
  assign _16545_ = \bapg_rd.w_ptr_r [2] ? _16544_ : _16541_;
  assign _16546_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[137] [15] : \MSYNC_1r1w.synth.nz.mem[136] [15];
  assign _16547_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[139] [15] : \MSYNC_1r1w.synth.nz.mem[138] [15];
  assign _16548_ = \bapg_rd.w_ptr_r [1] ? _16547_ : _16546_;
  assign _16549_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[141] [15] : \MSYNC_1r1w.synth.nz.mem[140] [15];
  assign _16550_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[143] [15] : \MSYNC_1r1w.synth.nz.mem[142] [15];
  assign _16551_ = \bapg_rd.w_ptr_r [1] ? _16550_ : _16549_;
  assign _16552_ = \bapg_rd.w_ptr_r [2] ? _16551_ : _16548_;
  assign _16553_ = \bapg_rd.w_ptr_r [3] ? _16552_ : _16545_;
  assign _16554_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[145] [15] : \MSYNC_1r1w.synth.nz.mem[144] [15];
  assign _16555_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[147] [15] : \MSYNC_1r1w.synth.nz.mem[146] [15];
  assign _16556_ = \bapg_rd.w_ptr_r [1] ? _16555_ : _16554_;
  assign _16557_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[149] [15] : \MSYNC_1r1w.synth.nz.mem[148] [15];
  assign _16558_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[151] [15] : \MSYNC_1r1w.synth.nz.mem[150] [15];
  assign _16559_ = \bapg_rd.w_ptr_r [1] ? _16558_ : _16557_;
  assign _16560_ = \bapg_rd.w_ptr_r [2] ? _16559_ : _16556_;
  assign _16561_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[153] [15] : \MSYNC_1r1w.synth.nz.mem[152] [15];
  assign _16562_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[155] [15] : \MSYNC_1r1w.synth.nz.mem[154] [15];
  assign _16563_ = \bapg_rd.w_ptr_r [1] ? _16562_ : _16561_;
  assign _16564_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[157] [15] : \MSYNC_1r1w.synth.nz.mem[156] [15];
  assign _16565_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[159] [15] : \MSYNC_1r1w.synth.nz.mem[158] [15];
  assign _16566_ = \bapg_rd.w_ptr_r [1] ? _16565_ : _16564_;
  assign _16567_ = \bapg_rd.w_ptr_r [2] ? _16566_ : _16563_;
  assign _16568_ = \bapg_rd.w_ptr_r [3] ? _16567_ : _16560_;
  assign _16569_ = \bapg_rd.w_ptr_r [4] ? _16568_ : _16553_;
  assign _16570_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[161] [15] : \MSYNC_1r1w.synth.nz.mem[160] [15];
  assign _16571_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[163] [15] : \MSYNC_1r1w.synth.nz.mem[162] [15];
  assign _16572_ = \bapg_rd.w_ptr_r [1] ? _16571_ : _16570_;
  assign _16573_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[165] [15] : \MSYNC_1r1w.synth.nz.mem[164] [15];
  assign _16574_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[167] [15] : \MSYNC_1r1w.synth.nz.mem[166] [15];
  assign _16575_ = \bapg_rd.w_ptr_r [1] ? _16574_ : _16573_;
  assign _16576_ = \bapg_rd.w_ptr_r [2] ? _16575_ : _16572_;
  assign _16577_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[169] [15] : \MSYNC_1r1w.synth.nz.mem[168] [15];
  assign _16578_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[171] [15] : \MSYNC_1r1w.synth.nz.mem[170] [15];
  assign _16579_ = \bapg_rd.w_ptr_r [1] ? _16578_ : _16577_;
  assign _16580_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[173] [15] : \MSYNC_1r1w.synth.nz.mem[172] [15];
  assign _16581_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[175] [15] : \MSYNC_1r1w.synth.nz.mem[174] [15];
  assign _16582_ = \bapg_rd.w_ptr_r [1] ? _16581_ : _16580_;
  assign _16583_ = \bapg_rd.w_ptr_r [2] ? _16582_ : _16579_;
  assign _16584_ = \bapg_rd.w_ptr_r [3] ? _16583_ : _16576_;
  assign _16585_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[177] [15] : \MSYNC_1r1w.synth.nz.mem[176] [15];
  assign _16586_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[179] [15] : \MSYNC_1r1w.synth.nz.mem[178] [15];
  assign _16587_ = \bapg_rd.w_ptr_r [1] ? _16586_ : _16585_;
  assign _16588_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[181] [15] : \MSYNC_1r1w.synth.nz.mem[180] [15];
  assign _16589_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[183] [15] : \MSYNC_1r1w.synth.nz.mem[182] [15];
  assign _16590_ = \bapg_rd.w_ptr_r [1] ? _16589_ : _16588_;
  assign _16591_ = \bapg_rd.w_ptr_r [2] ? _16590_ : _16587_;
  assign _16592_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[185] [15] : \MSYNC_1r1w.synth.nz.mem[184] [15];
  assign _16593_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[187] [15] : \MSYNC_1r1w.synth.nz.mem[186] [15];
  assign _16594_ = \bapg_rd.w_ptr_r [1] ? _16593_ : _16592_;
  assign _16595_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[189] [15] : \MSYNC_1r1w.synth.nz.mem[188] [15];
  assign _16596_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[191] [15] : \MSYNC_1r1w.synth.nz.mem[190] [15];
  assign _16597_ = \bapg_rd.w_ptr_r [1] ? _16596_ : _16595_;
  assign _16598_ = \bapg_rd.w_ptr_r [2] ? _16597_ : _16594_;
  assign _16599_ = \bapg_rd.w_ptr_r [3] ? _16598_ : _16591_;
  assign _16600_ = \bapg_rd.w_ptr_r [4] ? _16599_ : _16584_;
  assign _16601_ = \bapg_rd.w_ptr_r [5] ? _16600_ : _16569_;
  assign _16602_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[193] [15] : \MSYNC_1r1w.synth.nz.mem[192] [15];
  assign _16603_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[195] [15] : \MSYNC_1r1w.synth.nz.mem[194] [15];
  assign _16604_ = \bapg_rd.w_ptr_r [1] ? _16603_ : _16602_;
  assign _16605_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[197] [15] : \MSYNC_1r1w.synth.nz.mem[196] [15];
  assign _16606_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[199] [15] : \MSYNC_1r1w.synth.nz.mem[198] [15];
  assign _16607_ = \bapg_rd.w_ptr_r [1] ? _16606_ : _16605_;
  assign _16608_ = \bapg_rd.w_ptr_r [2] ? _16607_ : _16604_;
  assign _16609_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[201] [15] : \MSYNC_1r1w.synth.nz.mem[200] [15];
  assign _16610_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[203] [15] : \MSYNC_1r1w.synth.nz.mem[202] [15];
  assign _16611_ = \bapg_rd.w_ptr_r [1] ? _16610_ : _16609_;
  assign _16612_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[205] [15] : \MSYNC_1r1w.synth.nz.mem[204] [15];
  assign _16613_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[207] [15] : \MSYNC_1r1w.synth.nz.mem[206] [15];
  assign _16614_ = \bapg_rd.w_ptr_r [1] ? _16613_ : _16612_;
  assign _16615_ = \bapg_rd.w_ptr_r [2] ? _16614_ : _16611_;
  assign _16616_ = \bapg_rd.w_ptr_r [3] ? _16615_ : _16608_;
  assign _16617_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[209] [15] : \MSYNC_1r1w.synth.nz.mem[208] [15];
  assign _16618_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[211] [15] : \MSYNC_1r1w.synth.nz.mem[210] [15];
  assign _16619_ = \bapg_rd.w_ptr_r [1] ? _16618_ : _16617_;
  assign _16620_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[213] [15] : \MSYNC_1r1w.synth.nz.mem[212] [15];
  assign _16621_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[215] [15] : \MSYNC_1r1w.synth.nz.mem[214] [15];
  assign _16622_ = \bapg_rd.w_ptr_r [1] ? _16621_ : _16620_;
  assign _16623_ = \bapg_rd.w_ptr_r [2] ? _16622_ : _16619_;
  assign _16624_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[217] [15] : \MSYNC_1r1w.synth.nz.mem[216] [15];
  assign _16625_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[219] [15] : \MSYNC_1r1w.synth.nz.mem[218] [15];
  assign _16626_ = \bapg_rd.w_ptr_r [1] ? _16625_ : _16624_;
  assign _16627_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[221] [15] : \MSYNC_1r1w.synth.nz.mem[220] [15];
  assign _16628_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[223] [15] : \MSYNC_1r1w.synth.nz.mem[222] [15];
  assign _16629_ = \bapg_rd.w_ptr_r [1] ? _16628_ : _16627_;
  assign _16630_ = \bapg_rd.w_ptr_r [2] ? _16629_ : _16626_;
  assign _16631_ = \bapg_rd.w_ptr_r [3] ? _16630_ : _16623_;
  assign _16632_ = \bapg_rd.w_ptr_r [4] ? _16631_ : _16616_;
  assign _16633_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[225] [15] : \MSYNC_1r1w.synth.nz.mem[224] [15];
  assign _16634_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[227] [15] : \MSYNC_1r1w.synth.nz.mem[226] [15];
  assign _16635_ = \bapg_rd.w_ptr_r [1] ? _16634_ : _16633_;
  assign _16636_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[229] [15] : \MSYNC_1r1w.synth.nz.mem[228] [15];
  assign _16637_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[231] [15] : \MSYNC_1r1w.synth.nz.mem[230] [15];
  assign _16638_ = \bapg_rd.w_ptr_r [1] ? _16637_ : _16636_;
  assign _16639_ = \bapg_rd.w_ptr_r [2] ? _16638_ : _16635_;
  assign _16640_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[233] [15] : \MSYNC_1r1w.synth.nz.mem[232] [15];
  assign _16641_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[235] [15] : \MSYNC_1r1w.synth.nz.mem[234] [15];
  assign _16642_ = \bapg_rd.w_ptr_r [1] ? _16641_ : _16640_;
  assign _16643_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[237] [15] : \MSYNC_1r1w.synth.nz.mem[236] [15];
  assign _16644_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[239] [15] : \MSYNC_1r1w.synth.nz.mem[238] [15];
  assign _16645_ = \bapg_rd.w_ptr_r [1] ? _16644_ : _16643_;
  assign _16646_ = \bapg_rd.w_ptr_r [2] ? _16645_ : _16642_;
  assign _16647_ = \bapg_rd.w_ptr_r [3] ? _16646_ : _16639_;
  assign _16648_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[241] [15] : \MSYNC_1r1w.synth.nz.mem[240] [15];
  assign _16649_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[243] [15] : \MSYNC_1r1w.synth.nz.mem[242] [15];
  assign _16650_ = \bapg_rd.w_ptr_r [1] ? _16649_ : _16648_;
  assign _16651_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[245] [15] : \MSYNC_1r1w.synth.nz.mem[244] [15];
  assign _16652_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[247] [15] : \MSYNC_1r1w.synth.nz.mem[246] [15];
  assign _16653_ = \bapg_rd.w_ptr_r [1] ? _16652_ : _16651_;
  assign _16654_ = \bapg_rd.w_ptr_r [2] ? _16653_ : _16650_;
  assign _16655_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[249] [15] : \MSYNC_1r1w.synth.nz.mem[248] [15];
  assign _16656_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[251] [15] : \MSYNC_1r1w.synth.nz.mem[250] [15];
  assign _16657_ = \bapg_rd.w_ptr_r [1] ? _16656_ : _16655_;
  assign _16658_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[253] [15] : \MSYNC_1r1w.synth.nz.mem[252] [15];
  assign _16659_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[255] [15] : \MSYNC_1r1w.synth.nz.mem[254] [15];
  assign _16660_ = \bapg_rd.w_ptr_r [1] ? _16659_ : _16658_;
  assign _16661_ = \bapg_rd.w_ptr_r [2] ? _16660_ : _16657_;
  assign _16662_ = \bapg_rd.w_ptr_r [3] ? _16661_ : _16654_;
  assign _16663_ = \bapg_rd.w_ptr_r [4] ? _16662_ : _16647_;
  assign _16664_ = \bapg_rd.w_ptr_r [5] ? _16663_ : _16632_;
  assign _16665_ = \bapg_rd.w_ptr_r [6] ? _16664_ : _16601_;
  assign _16666_ = \bapg_rd.w_ptr_r [7] ? _16665_ : _16538_;
  assign _16667_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[257] [15] : \MSYNC_1r1w.synth.nz.mem[256] [15];
  assign _16668_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[259] [15] : \MSYNC_1r1w.synth.nz.mem[258] [15];
  assign _16669_ = \bapg_rd.w_ptr_r [1] ? _16668_ : _16667_;
  assign _16670_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[261] [15] : \MSYNC_1r1w.synth.nz.mem[260] [15];
  assign _16671_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[263] [15] : \MSYNC_1r1w.synth.nz.mem[262] [15];
  assign _16672_ = \bapg_rd.w_ptr_r [1] ? _16671_ : _16670_;
  assign _16673_ = \bapg_rd.w_ptr_r [2] ? _16672_ : _16669_;
  assign _16674_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[265] [15] : \MSYNC_1r1w.synth.nz.mem[264] [15];
  assign _16675_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[267] [15] : \MSYNC_1r1w.synth.nz.mem[266] [15];
  assign _16676_ = \bapg_rd.w_ptr_r [1] ? _16675_ : _16674_;
  assign _16677_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[269] [15] : \MSYNC_1r1w.synth.nz.mem[268] [15];
  assign _16678_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[271] [15] : \MSYNC_1r1w.synth.nz.mem[270] [15];
  assign _16679_ = \bapg_rd.w_ptr_r [1] ? _16678_ : _16677_;
  assign _16680_ = \bapg_rd.w_ptr_r [2] ? _16679_ : _16676_;
  assign _16681_ = \bapg_rd.w_ptr_r [3] ? _16680_ : _16673_;
  assign _16682_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[273] [15] : \MSYNC_1r1w.synth.nz.mem[272] [15];
  assign _16683_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[275] [15] : \MSYNC_1r1w.synth.nz.mem[274] [15];
  assign _16684_ = \bapg_rd.w_ptr_r [1] ? _16683_ : _16682_;
  assign _16685_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[277] [15] : \MSYNC_1r1w.synth.nz.mem[276] [15];
  assign _16686_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[279] [15] : \MSYNC_1r1w.synth.nz.mem[278] [15];
  assign _16687_ = \bapg_rd.w_ptr_r [1] ? _16686_ : _16685_;
  assign _16688_ = \bapg_rd.w_ptr_r [2] ? _16687_ : _16684_;
  assign _16689_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[281] [15] : \MSYNC_1r1w.synth.nz.mem[280] [15];
  assign _16690_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[283] [15] : \MSYNC_1r1w.synth.nz.mem[282] [15];
  assign _16691_ = \bapg_rd.w_ptr_r [1] ? _16690_ : _16689_;
  assign _16692_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[285] [15] : \MSYNC_1r1w.synth.nz.mem[284] [15];
  assign _16693_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[287] [15] : \MSYNC_1r1w.synth.nz.mem[286] [15];
  assign _16694_ = \bapg_rd.w_ptr_r [1] ? _16693_ : _16692_;
  assign _16695_ = \bapg_rd.w_ptr_r [2] ? _16694_ : _16691_;
  assign _16696_ = \bapg_rd.w_ptr_r [3] ? _16695_ : _16688_;
  assign _16697_ = \bapg_rd.w_ptr_r [4] ? _16696_ : _16681_;
  assign _16698_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[289] [15] : \MSYNC_1r1w.synth.nz.mem[288] [15];
  assign _16699_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[291] [15] : \MSYNC_1r1w.synth.nz.mem[290] [15];
  assign _16700_ = \bapg_rd.w_ptr_r [1] ? _16699_ : _16698_;
  assign _16701_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[293] [15] : \MSYNC_1r1w.synth.nz.mem[292] [15];
  assign _16702_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[295] [15] : \MSYNC_1r1w.synth.nz.mem[294] [15];
  assign _16703_ = \bapg_rd.w_ptr_r [1] ? _16702_ : _16701_;
  assign _16704_ = \bapg_rd.w_ptr_r [2] ? _16703_ : _16700_;
  assign _16705_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[297] [15] : \MSYNC_1r1w.synth.nz.mem[296] [15];
  assign _16706_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[299] [15] : \MSYNC_1r1w.synth.nz.mem[298] [15];
  assign _16707_ = \bapg_rd.w_ptr_r [1] ? _16706_ : _16705_;
  assign _16708_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[301] [15] : \MSYNC_1r1w.synth.nz.mem[300] [15];
  assign _16709_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[303] [15] : \MSYNC_1r1w.synth.nz.mem[302] [15];
  assign _16710_ = \bapg_rd.w_ptr_r [1] ? _16709_ : _16708_;
  assign _16711_ = \bapg_rd.w_ptr_r [2] ? _16710_ : _16707_;
  assign _16712_ = \bapg_rd.w_ptr_r [3] ? _16711_ : _16704_;
  assign _16713_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[305] [15] : \MSYNC_1r1w.synth.nz.mem[304] [15];
  assign _16714_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[307] [15] : \MSYNC_1r1w.synth.nz.mem[306] [15];
  assign _16715_ = \bapg_rd.w_ptr_r [1] ? _16714_ : _16713_;
  assign _16716_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[309] [15] : \MSYNC_1r1w.synth.nz.mem[308] [15];
  assign _16717_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[311] [15] : \MSYNC_1r1w.synth.nz.mem[310] [15];
  assign _16718_ = \bapg_rd.w_ptr_r [1] ? _16717_ : _16716_;
  assign _16719_ = \bapg_rd.w_ptr_r [2] ? _16718_ : _16715_;
  assign _16720_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[313] [15] : \MSYNC_1r1w.synth.nz.mem[312] [15];
  assign _16721_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[315] [15] : \MSYNC_1r1w.synth.nz.mem[314] [15];
  assign _16722_ = \bapg_rd.w_ptr_r [1] ? _16721_ : _16720_;
  assign _16723_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[317] [15] : \MSYNC_1r1w.synth.nz.mem[316] [15];
  assign _16724_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[319] [15] : \MSYNC_1r1w.synth.nz.mem[318] [15];
  assign _16725_ = \bapg_rd.w_ptr_r [1] ? _16724_ : _16723_;
  assign _16726_ = \bapg_rd.w_ptr_r [2] ? _16725_ : _16722_;
  assign _16727_ = \bapg_rd.w_ptr_r [3] ? _16726_ : _16719_;
  assign _16728_ = \bapg_rd.w_ptr_r [4] ? _16727_ : _16712_;
  assign _16729_ = \bapg_rd.w_ptr_r [5] ? _16728_ : _16697_;
  assign _16730_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[321] [15] : \MSYNC_1r1w.synth.nz.mem[320] [15];
  assign _16731_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[323] [15] : \MSYNC_1r1w.synth.nz.mem[322] [15];
  assign _16732_ = \bapg_rd.w_ptr_r [1] ? _16731_ : _16730_;
  assign _16733_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[325] [15] : \MSYNC_1r1w.synth.nz.mem[324] [15];
  assign _16734_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[327] [15] : \MSYNC_1r1w.synth.nz.mem[326] [15];
  assign _16735_ = \bapg_rd.w_ptr_r [1] ? _16734_ : _16733_;
  assign _16736_ = \bapg_rd.w_ptr_r [2] ? _16735_ : _16732_;
  assign _16737_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[329] [15] : \MSYNC_1r1w.synth.nz.mem[328] [15];
  assign _16738_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[331] [15] : \MSYNC_1r1w.synth.nz.mem[330] [15];
  assign _16739_ = \bapg_rd.w_ptr_r [1] ? _16738_ : _16737_;
  assign _16740_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[333] [15] : \MSYNC_1r1w.synth.nz.mem[332] [15];
  assign _16741_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[335] [15] : \MSYNC_1r1w.synth.nz.mem[334] [15];
  assign _16742_ = \bapg_rd.w_ptr_r [1] ? _16741_ : _16740_;
  assign _16743_ = \bapg_rd.w_ptr_r [2] ? _16742_ : _16739_;
  assign _16744_ = \bapg_rd.w_ptr_r [3] ? _16743_ : _16736_;
  assign _16745_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[337] [15] : \MSYNC_1r1w.synth.nz.mem[336] [15];
  assign _16746_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[339] [15] : \MSYNC_1r1w.synth.nz.mem[338] [15];
  assign _16747_ = \bapg_rd.w_ptr_r [1] ? _16746_ : _16745_;
  assign _16748_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[341] [15] : \MSYNC_1r1w.synth.nz.mem[340] [15];
  assign _16749_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[343] [15] : \MSYNC_1r1w.synth.nz.mem[342] [15];
  assign _16750_ = \bapg_rd.w_ptr_r [1] ? _16749_ : _16748_;
  assign _16751_ = \bapg_rd.w_ptr_r [2] ? _16750_ : _16747_;
  assign _16752_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[345] [15] : \MSYNC_1r1w.synth.nz.mem[344] [15];
  assign _16753_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[347] [15] : \MSYNC_1r1w.synth.nz.mem[346] [15];
  assign _16754_ = \bapg_rd.w_ptr_r [1] ? _16753_ : _16752_;
  assign _16755_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[349] [15] : \MSYNC_1r1w.synth.nz.mem[348] [15];
  assign _16756_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[351] [15] : \MSYNC_1r1w.synth.nz.mem[350] [15];
  assign _16757_ = \bapg_rd.w_ptr_r [1] ? _16756_ : _16755_;
  assign _16758_ = \bapg_rd.w_ptr_r [2] ? _16757_ : _16754_;
  assign _16759_ = \bapg_rd.w_ptr_r [3] ? _16758_ : _16751_;
  assign _16760_ = \bapg_rd.w_ptr_r [4] ? _16759_ : _16744_;
  assign _16761_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[353] [15] : \MSYNC_1r1w.synth.nz.mem[352] [15];
  assign _16762_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[355] [15] : \MSYNC_1r1w.synth.nz.mem[354] [15];
  assign _16763_ = \bapg_rd.w_ptr_r [1] ? _16762_ : _16761_;
  assign _16764_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[357] [15] : \MSYNC_1r1w.synth.nz.mem[356] [15];
  assign _16765_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[359] [15] : \MSYNC_1r1w.synth.nz.mem[358] [15];
  assign _16766_ = \bapg_rd.w_ptr_r [1] ? _16765_ : _16764_;
  assign _16767_ = \bapg_rd.w_ptr_r [2] ? _16766_ : _16763_;
  assign _16768_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[361] [15] : \MSYNC_1r1w.synth.nz.mem[360] [15];
  assign _16769_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[363] [15] : \MSYNC_1r1w.synth.nz.mem[362] [15];
  assign _16770_ = \bapg_rd.w_ptr_r [1] ? _16769_ : _16768_;
  assign _16771_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[365] [15] : \MSYNC_1r1w.synth.nz.mem[364] [15];
  assign _16772_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[367] [15] : \MSYNC_1r1w.synth.nz.mem[366] [15];
  assign _16773_ = \bapg_rd.w_ptr_r [1] ? _16772_ : _16771_;
  assign _16774_ = \bapg_rd.w_ptr_r [2] ? _16773_ : _16770_;
  assign _16775_ = \bapg_rd.w_ptr_r [3] ? _16774_ : _16767_;
  assign _16776_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[369] [15] : \MSYNC_1r1w.synth.nz.mem[368] [15];
  assign _16777_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[371] [15] : \MSYNC_1r1w.synth.nz.mem[370] [15];
  assign _16778_ = \bapg_rd.w_ptr_r [1] ? _16777_ : _16776_;
  assign _16779_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[373] [15] : \MSYNC_1r1w.synth.nz.mem[372] [15];
  assign _16780_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[375] [15] : \MSYNC_1r1w.synth.nz.mem[374] [15];
  assign _16781_ = \bapg_rd.w_ptr_r [1] ? _16780_ : _16779_;
  assign _16782_ = \bapg_rd.w_ptr_r [2] ? _16781_ : _16778_;
  assign _16783_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[377] [15] : \MSYNC_1r1w.synth.nz.mem[376] [15];
  assign _16784_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[379] [15] : \MSYNC_1r1w.synth.nz.mem[378] [15];
  assign _16785_ = \bapg_rd.w_ptr_r [1] ? _16784_ : _16783_;
  assign _16786_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[381] [15] : \MSYNC_1r1w.synth.nz.mem[380] [15];
  assign _16787_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[383] [15] : \MSYNC_1r1w.synth.nz.mem[382] [15];
  assign _16788_ = \bapg_rd.w_ptr_r [1] ? _16787_ : _16786_;
  assign _16789_ = \bapg_rd.w_ptr_r [2] ? _16788_ : _16785_;
  assign _16790_ = \bapg_rd.w_ptr_r [3] ? _16789_ : _16782_;
  assign _16791_ = \bapg_rd.w_ptr_r [4] ? _16790_ : _16775_;
  assign _16792_ = \bapg_rd.w_ptr_r [5] ? _16791_ : _16760_;
  assign _16793_ = \bapg_rd.w_ptr_r [6] ? _16792_ : _16729_;
  assign _16794_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[385] [15] : \MSYNC_1r1w.synth.nz.mem[384] [15];
  assign _16795_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[387] [15] : \MSYNC_1r1w.synth.nz.mem[386] [15];
  assign _16796_ = \bapg_rd.w_ptr_r [1] ? _16795_ : _16794_;
  assign _16797_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[389] [15] : \MSYNC_1r1w.synth.nz.mem[388] [15];
  assign _16798_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[391] [15] : \MSYNC_1r1w.synth.nz.mem[390] [15];
  assign _16799_ = \bapg_rd.w_ptr_r [1] ? _16798_ : _16797_;
  assign _16800_ = \bapg_rd.w_ptr_r [2] ? _16799_ : _16796_;
  assign _16801_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[393] [15] : \MSYNC_1r1w.synth.nz.mem[392] [15];
  assign _16802_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[395] [15] : \MSYNC_1r1w.synth.nz.mem[394] [15];
  assign _16803_ = \bapg_rd.w_ptr_r [1] ? _16802_ : _16801_;
  assign _16804_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[397] [15] : \MSYNC_1r1w.synth.nz.mem[396] [15];
  assign _16805_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[399] [15] : \MSYNC_1r1w.synth.nz.mem[398] [15];
  assign _16806_ = \bapg_rd.w_ptr_r [1] ? _16805_ : _16804_;
  assign _16807_ = \bapg_rd.w_ptr_r [2] ? _16806_ : _16803_;
  assign _16808_ = \bapg_rd.w_ptr_r [3] ? _16807_ : _16800_;
  assign _16809_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[401] [15] : \MSYNC_1r1w.synth.nz.mem[400] [15];
  assign _16810_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[403] [15] : \MSYNC_1r1w.synth.nz.mem[402] [15];
  assign _16811_ = \bapg_rd.w_ptr_r [1] ? _16810_ : _16809_;
  assign _16812_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[405] [15] : \MSYNC_1r1w.synth.nz.mem[404] [15];
  assign _16813_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[407] [15] : \MSYNC_1r1w.synth.nz.mem[406] [15];
  assign _16814_ = \bapg_rd.w_ptr_r [1] ? _16813_ : _16812_;
  assign _16815_ = \bapg_rd.w_ptr_r [2] ? _16814_ : _16811_;
  assign _16816_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[409] [15] : \MSYNC_1r1w.synth.nz.mem[408] [15];
  assign _16817_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[411] [15] : \MSYNC_1r1w.synth.nz.mem[410] [15];
  assign _16818_ = \bapg_rd.w_ptr_r [1] ? _16817_ : _16816_;
  assign _16819_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[413] [15] : \MSYNC_1r1w.synth.nz.mem[412] [15];
  assign _16820_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[415] [15] : \MSYNC_1r1w.synth.nz.mem[414] [15];
  assign _16821_ = \bapg_rd.w_ptr_r [1] ? _16820_ : _16819_;
  assign _16822_ = \bapg_rd.w_ptr_r [2] ? _16821_ : _16818_;
  assign _16823_ = \bapg_rd.w_ptr_r [3] ? _16822_ : _16815_;
  assign _16824_ = \bapg_rd.w_ptr_r [4] ? _16823_ : _16808_;
  assign _16825_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[417] [15] : \MSYNC_1r1w.synth.nz.mem[416] [15];
  assign _16826_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[419] [15] : \MSYNC_1r1w.synth.nz.mem[418] [15];
  assign _16827_ = \bapg_rd.w_ptr_r [1] ? _16826_ : _16825_;
  assign _16828_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[421] [15] : \MSYNC_1r1w.synth.nz.mem[420] [15];
  assign _16829_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[423] [15] : \MSYNC_1r1w.synth.nz.mem[422] [15];
  assign _16830_ = \bapg_rd.w_ptr_r [1] ? _16829_ : _16828_;
  assign _16831_ = \bapg_rd.w_ptr_r [2] ? _16830_ : _16827_;
  assign _16832_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[425] [15] : \MSYNC_1r1w.synth.nz.mem[424] [15];
  assign _16833_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[427] [15] : \MSYNC_1r1w.synth.nz.mem[426] [15];
  assign _16834_ = \bapg_rd.w_ptr_r [1] ? _16833_ : _16832_;
  assign _16835_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[429] [15] : \MSYNC_1r1w.synth.nz.mem[428] [15];
  assign _16836_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[431] [15] : \MSYNC_1r1w.synth.nz.mem[430] [15];
  assign _16837_ = \bapg_rd.w_ptr_r [1] ? _16836_ : _16835_;
  assign _16838_ = \bapg_rd.w_ptr_r [2] ? _16837_ : _16834_;
  assign _16839_ = \bapg_rd.w_ptr_r [3] ? _16838_ : _16831_;
  assign _16840_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[433] [15] : \MSYNC_1r1w.synth.nz.mem[432] [15];
  assign _16841_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[435] [15] : \MSYNC_1r1w.synth.nz.mem[434] [15];
  assign _16842_ = \bapg_rd.w_ptr_r [1] ? _16841_ : _16840_;
  assign _16843_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[437] [15] : \MSYNC_1r1w.synth.nz.mem[436] [15];
  assign _16844_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[439] [15] : \MSYNC_1r1w.synth.nz.mem[438] [15];
  assign _16845_ = \bapg_rd.w_ptr_r [1] ? _16844_ : _16843_;
  assign _16846_ = \bapg_rd.w_ptr_r [2] ? _16845_ : _16842_;
  assign _16847_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[441] [15] : \MSYNC_1r1w.synth.nz.mem[440] [15];
  assign _16848_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[443] [15] : \MSYNC_1r1w.synth.nz.mem[442] [15];
  assign _16849_ = \bapg_rd.w_ptr_r [1] ? _16848_ : _16847_;
  assign _16850_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[445] [15] : \MSYNC_1r1w.synth.nz.mem[444] [15];
  assign _16851_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[447] [15] : \MSYNC_1r1w.synth.nz.mem[446] [15];
  assign _16852_ = \bapg_rd.w_ptr_r [1] ? _16851_ : _16850_;
  assign _16853_ = \bapg_rd.w_ptr_r [2] ? _16852_ : _16849_;
  assign _16854_ = \bapg_rd.w_ptr_r [3] ? _16853_ : _16846_;
  assign _16855_ = \bapg_rd.w_ptr_r [4] ? _16854_ : _16839_;
  assign _16856_ = \bapg_rd.w_ptr_r [5] ? _16855_ : _16824_;
  assign _16857_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[449] [15] : \MSYNC_1r1w.synth.nz.mem[448] [15];
  assign _16858_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[451] [15] : \MSYNC_1r1w.synth.nz.mem[450] [15];
  assign _16859_ = \bapg_rd.w_ptr_r [1] ? _16858_ : _16857_;
  assign _16860_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[453] [15] : \MSYNC_1r1w.synth.nz.mem[452] [15];
  assign _16861_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[455] [15] : \MSYNC_1r1w.synth.nz.mem[454] [15];
  assign _16862_ = \bapg_rd.w_ptr_r [1] ? _16861_ : _16860_;
  assign _16863_ = \bapg_rd.w_ptr_r [2] ? _16862_ : _16859_;
  assign _16864_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[457] [15] : \MSYNC_1r1w.synth.nz.mem[456] [15];
  assign _16865_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[459] [15] : \MSYNC_1r1w.synth.nz.mem[458] [15];
  assign _16866_ = \bapg_rd.w_ptr_r [1] ? _16865_ : _16864_;
  assign _16867_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[461] [15] : \MSYNC_1r1w.synth.nz.mem[460] [15];
  assign _16868_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[463] [15] : \MSYNC_1r1w.synth.nz.mem[462] [15];
  assign _16869_ = \bapg_rd.w_ptr_r [1] ? _16868_ : _16867_;
  assign _16870_ = \bapg_rd.w_ptr_r [2] ? _16869_ : _16866_;
  assign _16871_ = \bapg_rd.w_ptr_r [3] ? _16870_ : _16863_;
  assign _16872_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[465] [15] : \MSYNC_1r1w.synth.nz.mem[464] [15];
  assign _16873_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[467] [15] : \MSYNC_1r1w.synth.nz.mem[466] [15];
  assign _16874_ = \bapg_rd.w_ptr_r [1] ? _16873_ : _16872_;
  assign _16875_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[469] [15] : \MSYNC_1r1w.synth.nz.mem[468] [15];
  assign _16876_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[471] [15] : \MSYNC_1r1w.synth.nz.mem[470] [15];
  assign _16877_ = \bapg_rd.w_ptr_r [1] ? _16876_ : _16875_;
  assign _16878_ = \bapg_rd.w_ptr_r [2] ? _16877_ : _16874_;
  assign _16879_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[473] [15] : \MSYNC_1r1w.synth.nz.mem[472] [15];
  assign _16880_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[475] [15] : \MSYNC_1r1w.synth.nz.mem[474] [15];
  assign _16881_ = \bapg_rd.w_ptr_r [1] ? _16880_ : _16879_;
  assign _16882_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[477] [15] : \MSYNC_1r1w.synth.nz.mem[476] [15];
  assign _16883_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[479] [15] : \MSYNC_1r1w.synth.nz.mem[478] [15];
  assign _16884_ = \bapg_rd.w_ptr_r [1] ? _16883_ : _16882_;
  assign _16885_ = \bapg_rd.w_ptr_r [2] ? _16884_ : _16881_;
  assign _16886_ = \bapg_rd.w_ptr_r [3] ? _16885_ : _16878_;
  assign _16887_ = \bapg_rd.w_ptr_r [4] ? _16886_ : _16871_;
  assign _16888_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[481] [15] : \MSYNC_1r1w.synth.nz.mem[480] [15];
  assign _16889_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[483] [15] : \MSYNC_1r1w.synth.nz.mem[482] [15];
  assign _16890_ = \bapg_rd.w_ptr_r [1] ? _16889_ : _16888_;
  assign _16891_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[485] [15] : \MSYNC_1r1w.synth.nz.mem[484] [15];
  assign _16892_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[487] [15] : \MSYNC_1r1w.synth.nz.mem[486] [15];
  assign _16893_ = \bapg_rd.w_ptr_r [1] ? _16892_ : _16891_;
  assign _16894_ = \bapg_rd.w_ptr_r [2] ? _16893_ : _16890_;
  assign _16895_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[489] [15] : \MSYNC_1r1w.synth.nz.mem[488] [15];
  assign _16896_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[491] [15] : \MSYNC_1r1w.synth.nz.mem[490] [15];
  assign _16897_ = \bapg_rd.w_ptr_r [1] ? _16896_ : _16895_;
  assign _16898_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[493] [15] : \MSYNC_1r1w.synth.nz.mem[492] [15];
  assign _16899_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[495] [15] : \MSYNC_1r1w.synth.nz.mem[494] [15];
  assign _16900_ = \bapg_rd.w_ptr_r [1] ? _16899_ : _16898_;
  assign _16901_ = \bapg_rd.w_ptr_r [2] ? _16900_ : _16897_;
  assign _16902_ = \bapg_rd.w_ptr_r [3] ? _16901_ : _16894_;
  assign _16903_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[497] [15] : \MSYNC_1r1w.synth.nz.mem[496] [15];
  assign _16904_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[499] [15] : \MSYNC_1r1w.synth.nz.mem[498] [15];
  assign _16905_ = \bapg_rd.w_ptr_r [1] ? _16904_ : _16903_;
  assign _16906_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[501] [15] : \MSYNC_1r1w.synth.nz.mem[500] [15];
  assign _16907_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[503] [15] : \MSYNC_1r1w.synth.nz.mem[502] [15];
  assign _16908_ = \bapg_rd.w_ptr_r [1] ? _16907_ : _16906_;
  assign _16909_ = \bapg_rd.w_ptr_r [2] ? _16908_ : _16905_;
  assign _16910_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[505] [15] : \MSYNC_1r1w.synth.nz.mem[504] [15];
  assign _16911_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[507] [15] : \MSYNC_1r1w.synth.nz.mem[506] [15];
  assign _16912_ = \bapg_rd.w_ptr_r [1] ? _16911_ : _16910_;
  assign _16913_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[509] [15] : \MSYNC_1r1w.synth.nz.mem[508] [15];
  assign _16914_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[511] [15] : \MSYNC_1r1w.synth.nz.mem[510] [15];
  assign _16915_ = \bapg_rd.w_ptr_r [1] ? _16914_ : _16913_;
  assign _16916_ = \bapg_rd.w_ptr_r [2] ? _16915_ : _16912_;
  assign _16917_ = \bapg_rd.w_ptr_r [3] ? _16916_ : _16909_;
  assign _16918_ = \bapg_rd.w_ptr_r [4] ? _16917_ : _16902_;
  assign _16919_ = \bapg_rd.w_ptr_r [5] ? _16918_ : _16887_;
  assign _16920_ = \bapg_rd.w_ptr_r [6] ? _16919_ : _16856_;
  assign _16921_ = \bapg_rd.w_ptr_r [7] ? _16920_ : _16793_;
  assign _16922_ = \bapg_rd.w_ptr_r [8] ? _16921_ : _16666_;
  assign _16923_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[513] [15] : \MSYNC_1r1w.synth.nz.mem[512] [15];
  assign _16924_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[515] [15] : \MSYNC_1r1w.synth.nz.mem[514] [15];
  assign _16925_ = \bapg_rd.w_ptr_r [1] ? _16924_ : _16923_;
  assign _16926_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[517] [15] : \MSYNC_1r1w.synth.nz.mem[516] [15];
  assign _16927_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[519] [15] : \MSYNC_1r1w.synth.nz.mem[518] [15];
  assign _16928_ = \bapg_rd.w_ptr_r [1] ? _16927_ : _16926_;
  assign _16929_ = \bapg_rd.w_ptr_r [2] ? _16928_ : _16925_;
  assign _16930_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[521] [15] : \MSYNC_1r1w.synth.nz.mem[520] [15];
  assign _16931_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[523] [15] : \MSYNC_1r1w.synth.nz.mem[522] [15];
  assign _16932_ = \bapg_rd.w_ptr_r [1] ? _16931_ : _16930_;
  assign _16933_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[525] [15] : \MSYNC_1r1w.synth.nz.mem[524] [15];
  assign _16934_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[527] [15] : \MSYNC_1r1w.synth.nz.mem[526] [15];
  assign _16935_ = \bapg_rd.w_ptr_r [1] ? _16934_ : _16933_;
  assign _16936_ = \bapg_rd.w_ptr_r [2] ? _16935_ : _16932_;
  assign _16937_ = \bapg_rd.w_ptr_r [3] ? _16936_ : _16929_;
  assign _16938_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[529] [15] : \MSYNC_1r1w.synth.nz.mem[528] [15];
  assign _16939_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[531] [15] : \MSYNC_1r1w.synth.nz.mem[530] [15];
  assign _16940_ = \bapg_rd.w_ptr_r [1] ? _16939_ : _16938_;
  assign _16941_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[533] [15] : \MSYNC_1r1w.synth.nz.mem[532] [15];
  assign _16942_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[535] [15] : \MSYNC_1r1w.synth.nz.mem[534] [15];
  assign _16943_ = \bapg_rd.w_ptr_r [1] ? _16942_ : _16941_;
  assign _16944_ = \bapg_rd.w_ptr_r [2] ? _16943_ : _16940_;
  assign _16945_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[537] [15] : \MSYNC_1r1w.synth.nz.mem[536] [15];
  assign _16946_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[539] [15] : \MSYNC_1r1w.synth.nz.mem[538] [15];
  assign _16947_ = \bapg_rd.w_ptr_r [1] ? _16946_ : _16945_;
  assign _16948_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[541] [15] : \MSYNC_1r1w.synth.nz.mem[540] [15];
  assign _16949_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[543] [15] : \MSYNC_1r1w.synth.nz.mem[542] [15];
  assign _16950_ = \bapg_rd.w_ptr_r [1] ? _16949_ : _16948_;
  assign _16951_ = \bapg_rd.w_ptr_r [2] ? _16950_ : _16947_;
  assign _16952_ = \bapg_rd.w_ptr_r [3] ? _16951_ : _16944_;
  assign _16953_ = \bapg_rd.w_ptr_r [4] ? _16952_ : _16937_;
  assign _16954_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[545] [15] : \MSYNC_1r1w.synth.nz.mem[544] [15];
  assign _16955_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[547] [15] : \MSYNC_1r1w.synth.nz.mem[546] [15];
  assign _16956_ = \bapg_rd.w_ptr_r [1] ? _16955_ : _16954_;
  assign _16957_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[549] [15] : \MSYNC_1r1w.synth.nz.mem[548] [15];
  assign _16958_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[551] [15] : \MSYNC_1r1w.synth.nz.mem[550] [15];
  assign _16959_ = \bapg_rd.w_ptr_r [1] ? _16958_ : _16957_;
  assign _16960_ = \bapg_rd.w_ptr_r [2] ? _16959_ : _16956_;
  assign _16961_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[553] [15] : \MSYNC_1r1w.synth.nz.mem[552] [15];
  assign _16962_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[555] [15] : \MSYNC_1r1w.synth.nz.mem[554] [15];
  assign _16963_ = \bapg_rd.w_ptr_r [1] ? _16962_ : _16961_;
  assign _16964_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[557] [15] : \MSYNC_1r1w.synth.nz.mem[556] [15];
  assign _16965_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[559] [15] : \MSYNC_1r1w.synth.nz.mem[558] [15];
  assign _16966_ = \bapg_rd.w_ptr_r [1] ? _16965_ : _16964_;
  assign _16967_ = \bapg_rd.w_ptr_r [2] ? _16966_ : _16963_;
  assign _16968_ = \bapg_rd.w_ptr_r [3] ? _16967_ : _16960_;
  assign _16969_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[561] [15] : \MSYNC_1r1w.synth.nz.mem[560] [15];
  assign _16970_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[563] [15] : \MSYNC_1r1w.synth.nz.mem[562] [15];
  assign _16971_ = \bapg_rd.w_ptr_r [1] ? _16970_ : _16969_;
  assign _16972_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[565] [15] : \MSYNC_1r1w.synth.nz.mem[564] [15];
  assign _16973_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[567] [15] : \MSYNC_1r1w.synth.nz.mem[566] [15];
  assign _16974_ = \bapg_rd.w_ptr_r [1] ? _16973_ : _16972_;
  assign _16975_ = \bapg_rd.w_ptr_r [2] ? _16974_ : _16971_;
  assign _16976_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[569] [15] : \MSYNC_1r1w.synth.nz.mem[568] [15];
  assign _16977_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[571] [15] : \MSYNC_1r1w.synth.nz.mem[570] [15];
  assign _16978_ = \bapg_rd.w_ptr_r [1] ? _16977_ : _16976_;
  assign _16979_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[573] [15] : \MSYNC_1r1w.synth.nz.mem[572] [15];
  assign _16980_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[575] [15] : \MSYNC_1r1w.synth.nz.mem[574] [15];
  assign _16981_ = \bapg_rd.w_ptr_r [1] ? _16980_ : _16979_;
  assign _16982_ = \bapg_rd.w_ptr_r [2] ? _16981_ : _16978_;
  assign _16983_ = \bapg_rd.w_ptr_r [3] ? _16982_ : _16975_;
  assign _16984_ = \bapg_rd.w_ptr_r [4] ? _16983_ : _16968_;
  assign _16985_ = \bapg_rd.w_ptr_r [5] ? _16984_ : _16953_;
  assign _16986_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[577] [15] : \MSYNC_1r1w.synth.nz.mem[576] [15];
  assign _16987_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[579] [15] : \MSYNC_1r1w.synth.nz.mem[578] [15];
  assign _16988_ = \bapg_rd.w_ptr_r [1] ? _16987_ : _16986_;
  assign _16989_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[581] [15] : \MSYNC_1r1w.synth.nz.mem[580] [15];
  assign _16990_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[583] [15] : \MSYNC_1r1w.synth.nz.mem[582] [15];
  assign _16991_ = \bapg_rd.w_ptr_r [1] ? _16990_ : _16989_;
  assign _16992_ = \bapg_rd.w_ptr_r [2] ? _16991_ : _16988_;
  assign _16993_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[585] [15] : \MSYNC_1r1w.synth.nz.mem[584] [15];
  assign _16994_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[587] [15] : \MSYNC_1r1w.synth.nz.mem[586] [15];
  assign _16995_ = \bapg_rd.w_ptr_r [1] ? _16994_ : _16993_;
  assign _16996_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[589] [15] : \MSYNC_1r1w.synth.nz.mem[588] [15];
  assign _16997_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[591] [15] : \MSYNC_1r1w.synth.nz.mem[590] [15];
  assign _16998_ = \bapg_rd.w_ptr_r [1] ? _16997_ : _16996_;
  assign _16999_ = \bapg_rd.w_ptr_r [2] ? _16998_ : _16995_;
  assign _17000_ = \bapg_rd.w_ptr_r [3] ? _16999_ : _16992_;
  assign _17001_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[593] [15] : \MSYNC_1r1w.synth.nz.mem[592] [15];
  assign _17002_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[595] [15] : \MSYNC_1r1w.synth.nz.mem[594] [15];
  assign _17003_ = \bapg_rd.w_ptr_r [1] ? _17002_ : _17001_;
  assign _17004_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[597] [15] : \MSYNC_1r1w.synth.nz.mem[596] [15];
  assign _17005_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[599] [15] : \MSYNC_1r1w.synth.nz.mem[598] [15];
  assign _17006_ = \bapg_rd.w_ptr_r [1] ? _17005_ : _17004_;
  assign _17007_ = \bapg_rd.w_ptr_r [2] ? _17006_ : _17003_;
  assign _17008_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[601] [15] : \MSYNC_1r1w.synth.nz.mem[600] [15];
  assign _17009_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[603] [15] : \MSYNC_1r1w.synth.nz.mem[602] [15];
  assign _17010_ = \bapg_rd.w_ptr_r [1] ? _17009_ : _17008_;
  assign _17011_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[605] [15] : \MSYNC_1r1w.synth.nz.mem[604] [15];
  assign _17012_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[607] [15] : \MSYNC_1r1w.synth.nz.mem[606] [15];
  assign _17013_ = \bapg_rd.w_ptr_r [1] ? _17012_ : _17011_;
  assign _17014_ = \bapg_rd.w_ptr_r [2] ? _17013_ : _17010_;
  assign _17015_ = \bapg_rd.w_ptr_r [3] ? _17014_ : _17007_;
  assign _17016_ = \bapg_rd.w_ptr_r [4] ? _17015_ : _17000_;
  assign _17017_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[609] [15] : \MSYNC_1r1w.synth.nz.mem[608] [15];
  assign _17018_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[611] [15] : \MSYNC_1r1w.synth.nz.mem[610] [15];
  assign _17019_ = \bapg_rd.w_ptr_r [1] ? _17018_ : _17017_;
  assign _17020_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[613] [15] : \MSYNC_1r1w.synth.nz.mem[612] [15];
  assign _17021_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[615] [15] : \MSYNC_1r1w.synth.nz.mem[614] [15];
  assign _17022_ = \bapg_rd.w_ptr_r [1] ? _17021_ : _17020_;
  assign _17023_ = \bapg_rd.w_ptr_r [2] ? _17022_ : _17019_;
  assign _17024_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[617] [15] : \MSYNC_1r1w.synth.nz.mem[616] [15];
  assign _17025_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[619] [15] : \MSYNC_1r1w.synth.nz.mem[618] [15];
  assign _17026_ = \bapg_rd.w_ptr_r [1] ? _17025_ : _17024_;
  assign _17027_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[621] [15] : \MSYNC_1r1w.synth.nz.mem[620] [15];
  assign _17028_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[623] [15] : \MSYNC_1r1w.synth.nz.mem[622] [15];
  assign _17029_ = \bapg_rd.w_ptr_r [1] ? _17028_ : _17027_;
  assign _17030_ = \bapg_rd.w_ptr_r [2] ? _17029_ : _17026_;
  assign _17031_ = \bapg_rd.w_ptr_r [3] ? _17030_ : _17023_;
  assign _17032_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[625] [15] : \MSYNC_1r1w.synth.nz.mem[624] [15];
  assign _17033_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[627] [15] : \MSYNC_1r1w.synth.nz.mem[626] [15];
  assign _17034_ = \bapg_rd.w_ptr_r [1] ? _17033_ : _17032_;
  assign _17035_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[629] [15] : \MSYNC_1r1w.synth.nz.mem[628] [15];
  assign _17036_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[631] [15] : \MSYNC_1r1w.synth.nz.mem[630] [15];
  assign _17037_ = \bapg_rd.w_ptr_r [1] ? _17036_ : _17035_;
  assign _17038_ = \bapg_rd.w_ptr_r [2] ? _17037_ : _17034_;
  assign _17039_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[633] [15] : \MSYNC_1r1w.synth.nz.mem[632] [15];
  assign _17040_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[635] [15] : \MSYNC_1r1w.synth.nz.mem[634] [15];
  assign _17041_ = \bapg_rd.w_ptr_r [1] ? _17040_ : _17039_;
  assign _17042_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[637] [15] : \MSYNC_1r1w.synth.nz.mem[636] [15];
  assign _17043_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[639] [15] : \MSYNC_1r1w.synth.nz.mem[638] [15];
  assign _17044_ = \bapg_rd.w_ptr_r [1] ? _17043_ : _17042_;
  assign _17045_ = \bapg_rd.w_ptr_r [2] ? _17044_ : _17041_;
  assign _17046_ = \bapg_rd.w_ptr_r [3] ? _17045_ : _17038_;
  assign _17047_ = \bapg_rd.w_ptr_r [4] ? _17046_ : _17031_;
  assign _17048_ = \bapg_rd.w_ptr_r [5] ? _17047_ : _17016_;
  assign _17049_ = \bapg_rd.w_ptr_r [6] ? _17048_ : _16985_;
  assign _17050_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[641] [15] : \MSYNC_1r1w.synth.nz.mem[640] [15];
  assign _17051_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[643] [15] : \MSYNC_1r1w.synth.nz.mem[642] [15];
  assign _17052_ = \bapg_rd.w_ptr_r [1] ? _17051_ : _17050_;
  assign _17053_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[645] [15] : \MSYNC_1r1w.synth.nz.mem[644] [15];
  assign _17054_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[647] [15] : \MSYNC_1r1w.synth.nz.mem[646] [15];
  assign _17055_ = \bapg_rd.w_ptr_r [1] ? _17054_ : _17053_;
  assign _17056_ = \bapg_rd.w_ptr_r [2] ? _17055_ : _17052_;
  assign _17057_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[649] [15] : \MSYNC_1r1w.synth.nz.mem[648] [15];
  assign _17058_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[651] [15] : \MSYNC_1r1w.synth.nz.mem[650] [15];
  assign _17059_ = \bapg_rd.w_ptr_r [1] ? _17058_ : _17057_;
  assign _17060_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[653] [15] : \MSYNC_1r1w.synth.nz.mem[652] [15];
  assign _17061_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[655] [15] : \MSYNC_1r1w.synth.nz.mem[654] [15];
  assign _17062_ = \bapg_rd.w_ptr_r [1] ? _17061_ : _17060_;
  assign _17063_ = \bapg_rd.w_ptr_r [2] ? _17062_ : _17059_;
  assign _17064_ = \bapg_rd.w_ptr_r [3] ? _17063_ : _17056_;
  assign _17065_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[657] [15] : \MSYNC_1r1w.synth.nz.mem[656] [15];
  assign _17066_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[659] [15] : \MSYNC_1r1w.synth.nz.mem[658] [15];
  assign _17067_ = \bapg_rd.w_ptr_r [1] ? _17066_ : _17065_;
  assign _17068_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[661] [15] : \MSYNC_1r1w.synth.nz.mem[660] [15];
  assign _17069_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[663] [15] : \MSYNC_1r1w.synth.nz.mem[662] [15];
  assign _17070_ = \bapg_rd.w_ptr_r [1] ? _17069_ : _17068_;
  assign _17071_ = \bapg_rd.w_ptr_r [2] ? _17070_ : _17067_;
  assign _17072_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[665] [15] : \MSYNC_1r1w.synth.nz.mem[664] [15];
  assign _17073_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[667] [15] : \MSYNC_1r1w.synth.nz.mem[666] [15];
  assign _17074_ = \bapg_rd.w_ptr_r [1] ? _17073_ : _17072_;
  assign _17075_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[669] [15] : \MSYNC_1r1w.synth.nz.mem[668] [15];
  assign _17076_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[671] [15] : \MSYNC_1r1w.synth.nz.mem[670] [15];
  assign _17077_ = \bapg_rd.w_ptr_r [1] ? _17076_ : _17075_;
  assign _17078_ = \bapg_rd.w_ptr_r [2] ? _17077_ : _17074_;
  assign _17079_ = \bapg_rd.w_ptr_r [3] ? _17078_ : _17071_;
  assign _17080_ = \bapg_rd.w_ptr_r [4] ? _17079_ : _17064_;
  assign _17081_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[673] [15] : \MSYNC_1r1w.synth.nz.mem[672] [15];
  assign _17082_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[675] [15] : \MSYNC_1r1w.synth.nz.mem[674] [15];
  assign _17083_ = \bapg_rd.w_ptr_r [1] ? _17082_ : _17081_;
  assign _17084_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[677] [15] : \MSYNC_1r1w.synth.nz.mem[676] [15];
  assign _17085_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[679] [15] : \MSYNC_1r1w.synth.nz.mem[678] [15];
  assign _17086_ = \bapg_rd.w_ptr_r [1] ? _17085_ : _17084_;
  assign _17087_ = \bapg_rd.w_ptr_r [2] ? _17086_ : _17083_;
  assign _17088_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[681] [15] : \MSYNC_1r1w.synth.nz.mem[680] [15];
  assign _17089_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[683] [15] : \MSYNC_1r1w.synth.nz.mem[682] [15];
  assign _17090_ = \bapg_rd.w_ptr_r [1] ? _17089_ : _17088_;
  assign _17091_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[685] [15] : \MSYNC_1r1w.synth.nz.mem[684] [15];
  assign _17092_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[687] [15] : \MSYNC_1r1w.synth.nz.mem[686] [15];
  assign _17093_ = \bapg_rd.w_ptr_r [1] ? _17092_ : _17091_;
  assign _17094_ = \bapg_rd.w_ptr_r [2] ? _17093_ : _17090_;
  assign _17095_ = \bapg_rd.w_ptr_r [3] ? _17094_ : _17087_;
  assign _17096_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[689] [15] : \MSYNC_1r1w.synth.nz.mem[688] [15];
  assign _17097_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[691] [15] : \MSYNC_1r1w.synth.nz.mem[690] [15];
  assign _17098_ = \bapg_rd.w_ptr_r [1] ? _17097_ : _17096_;
  assign _17099_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[693] [15] : \MSYNC_1r1w.synth.nz.mem[692] [15];
  assign _17100_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[695] [15] : \MSYNC_1r1w.synth.nz.mem[694] [15];
  assign _17101_ = \bapg_rd.w_ptr_r [1] ? _17100_ : _17099_;
  assign _17102_ = \bapg_rd.w_ptr_r [2] ? _17101_ : _17098_;
  assign _17103_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[697] [15] : \MSYNC_1r1w.synth.nz.mem[696] [15];
  assign _17104_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[699] [15] : \MSYNC_1r1w.synth.nz.mem[698] [15];
  assign _17105_ = \bapg_rd.w_ptr_r [1] ? _17104_ : _17103_;
  assign _17106_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[701] [15] : \MSYNC_1r1w.synth.nz.mem[700] [15];
  assign _17107_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[703] [15] : \MSYNC_1r1w.synth.nz.mem[702] [15];
  assign _17108_ = \bapg_rd.w_ptr_r [1] ? _17107_ : _17106_;
  assign _17109_ = \bapg_rd.w_ptr_r [2] ? _17108_ : _17105_;
  assign _17110_ = \bapg_rd.w_ptr_r [3] ? _17109_ : _17102_;
  assign _17111_ = \bapg_rd.w_ptr_r [4] ? _17110_ : _17095_;
  assign _17112_ = \bapg_rd.w_ptr_r [5] ? _17111_ : _17080_;
  assign _17113_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[705] [15] : \MSYNC_1r1w.synth.nz.mem[704] [15];
  assign _17114_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[707] [15] : \MSYNC_1r1w.synth.nz.mem[706] [15];
  assign _17115_ = \bapg_rd.w_ptr_r [1] ? _17114_ : _17113_;
  assign _17116_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[709] [15] : \MSYNC_1r1w.synth.nz.mem[708] [15];
  assign _17117_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[711] [15] : \MSYNC_1r1w.synth.nz.mem[710] [15];
  assign _17118_ = \bapg_rd.w_ptr_r [1] ? _17117_ : _17116_;
  assign _17119_ = \bapg_rd.w_ptr_r [2] ? _17118_ : _17115_;
  assign _17120_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[713] [15] : \MSYNC_1r1w.synth.nz.mem[712] [15];
  assign _17121_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[715] [15] : \MSYNC_1r1w.synth.nz.mem[714] [15];
  assign _17122_ = \bapg_rd.w_ptr_r [1] ? _17121_ : _17120_;
  assign _17123_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[717] [15] : \MSYNC_1r1w.synth.nz.mem[716] [15];
  assign _17124_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[719] [15] : \MSYNC_1r1w.synth.nz.mem[718] [15];
  assign _17125_ = \bapg_rd.w_ptr_r [1] ? _17124_ : _17123_;
  assign _17126_ = \bapg_rd.w_ptr_r [2] ? _17125_ : _17122_;
  assign _17127_ = \bapg_rd.w_ptr_r [3] ? _17126_ : _17119_;
  assign _17128_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[721] [15] : \MSYNC_1r1w.synth.nz.mem[720] [15];
  assign _17129_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[723] [15] : \MSYNC_1r1w.synth.nz.mem[722] [15];
  assign _17130_ = \bapg_rd.w_ptr_r [1] ? _17129_ : _17128_;
  assign _17131_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[725] [15] : \MSYNC_1r1w.synth.nz.mem[724] [15];
  assign _17132_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[727] [15] : \MSYNC_1r1w.synth.nz.mem[726] [15];
  assign _17133_ = \bapg_rd.w_ptr_r [1] ? _17132_ : _17131_;
  assign _17134_ = \bapg_rd.w_ptr_r [2] ? _17133_ : _17130_;
  assign _17135_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[729] [15] : \MSYNC_1r1w.synth.nz.mem[728] [15];
  assign _17136_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[731] [15] : \MSYNC_1r1w.synth.nz.mem[730] [15];
  assign _17137_ = \bapg_rd.w_ptr_r [1] ? _17136_ : _17135_;
  assign _17138_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[733] [15] : \MSYNC_1r1w.synth.nz.mem[732] [15];
  assign _17139_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[735] [15] : \MSYNC_1r1w.synth.nz.mem[734] [15];
  assign _17140_ = \bapg_rd.w_ptr_r [1] ? _17139_ : _17138_;
  assign _17141_ = \bapg_rd.w_ptr_r [2] ? _17140_ : _17137_;
  assign _17142_ = \bapg_rd.w_ptr_r [3] ? _17141_ : _17134_;
  assign _17143_ = \bapg_rd.w_ptr_r [4] ? _17142_ : _17127_;
  assign _17144_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[737] [15] : \MSYNC_1r1w.synth.nz.mem[736] [15];
  assign _17145_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[739] [15] : \MSYNC_1r1w.synth.nz.mem[738] [15];
  assign _17146_ = \bapg_rd.w_ptr_r [1] ? _17145_ : _17144_;
  assign _17147_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[741] [15] : \MSYNC_1r1w.synth.nz.mem[740] [15];
  assign _17148_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[743] [15] : \MSYNC_1r1w.synth.nz.mem[742] [15];
  assign _17149_ = \bapg_rd.w_ptr_r [1] ? _17148_ : _17147_;
  assign _17150_ = \bapg_rd.w_ptr_r [2] ? _17149_ : _17146_;
  assign _17151_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[745] [15] : \MSYNC_1r1w.synth.nz.mem[744] [15];
  assign _17152_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[747] [15] : \MSYNC_1r1w.synth.nz.mem[746] [15];
  assign _17153_ = \bapg_rd.w_ptr_r [1] ? _17152_ : _17151_;
  assign _17154_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[749] [15] : \MSYNC_1r1w.synth.nz.mem[748] [15];
  assign _17155_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[751] [15] : \MSYNC_1r1w.synth.nz.mem[750] [15];
  assign _17156_ = \bapg_rd.w_ptr_r [1] ? _17155_ : _17154_;
  assign _17157_ = \bapg_rd.w_ptr_r [2] ? _17156_ : _17153_;
  assign _17158_ = \bapg_rd.w_ptr_r [3] ? _17157_ : _17150_;
  assign _17159_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[753] [15] : \MSYNC_1r1w.synth.nz.mem[752] [15];
  assign _17160_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[755] [15] : \MSYNC_1r1w.synth.nz.mem[754] [15];
  assign _17161_ = \bapg_rd.w_ptr_r [1] ? _17160_ : _17159_;
  assign _17162_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[757] [15] : \MSYNC_1r1w.synth.nz.mem[756] [15];
  assign _17163_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[759] [15] : \MSYNC_1r1w.synth.nz.mem[758] [15];
  assign _17164_ = \bapg_rd.w_ptr_r [1] ? _17163_ : _17162_;
  assign _17165_ = \bapg_rd.w_ptr_r [2] ? _17164_ : _17161_;
  assign _17166_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[761] [15] : \MSYNC_1r1w.synth.nz.mem[760] [15];
  assign _17167_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[763] [15] : \MSYNC_1r1w.synth.nz.mem[762] [15];
  assign _17168_ = \bapg_rd.w_ptr_r [1] ? _17167_ : _17166_;
  assign _17169_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[765] [15] : \MSYNC_1r1w.synth.nz.mem[764] [15];
  assign _17170_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[767] [15] : \MSYNC_1r1w.synth.nz.mem[766] [15];
  assign _17171_ = \bapg_rd.w_ptr_r [1] ? _17170_ : _17169_;
  assign _17172_ = \bapg_rd.w_ptr_r [2] ? _17171_ : _17168_;
  assign _17173_ = \bapg_rd.w_ptr_r [3] ? _17172_ : _17165_;
  assign _17174_ = \bapg_rd.w_ptr_r [4] ? _17173_ : _17158_;
  assign _17175_ = \bapg_rd.w_ptr_r [5] ? _17174_ : _17143_;
  assign _17176_ = \bapg_rd.w_ptr_r [6] ? _17175_ : _17112_;
  assign _17177_ = \bapg_rd.w_ptr_r [7] ? _17176_ : _17049_;
  assign _17178_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[769] [15] : \MSYNC_1r1w.synth.nz.mem[768] [15];
  assign _17179_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[771] [15] : \MSYNC_1r1w.synth.nz.mem[770] [15];
  assign _17180_ = \bapg_rd.w_ptr_r [1] ? _17179_ : _17178_;
  assign _17181_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[773] [15] : \MSYNC_1r1w.synth.nz.mem[772] [15];
  assign _17182_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[775] [15] : \MSYNC_1r1w.synth.nz.mem[774] [15];
  assign _17183_ = \bapg_rd.w_ptr_r [1] ? _17182_ : _17181_;
  assign _17184_ = \bapg_rd.w_ptr_r [2] ? _17183_ : _17180_;
  assign _17185_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[777] [15] : \MSYNC_1r1w.synth.nz.mem[776] [15];
  assign _17186_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[779] [15] : \MSYNC_1r1w.synth.nz.mem[778] [15];
  assign _17187_ = \bapg_rd.w_ptr_r [1] ? _17186_ : _17185_;
  assign _17188_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[781] [15] : \MSYNC_1r1w.synth.nz.mem[780] [15];
  assign _17189_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[783] [15] : \MSYNC_1r1w.synth.nz.mem[782] [15];
  assign _17190_ = \bapg_rd.w_ptr_r [1] ? _17189_ : _17188_;
  assign _17191_ = \bapg_rd.w_ptr_r [2] ? _17190_ : _17187_;
  assign _17192_ = \bapg_rd.w_ptr_r [3] ? _17191_ : _17184_;
  assign _17193_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[785] [15] : \MSYNC_1r1w.synth.nz.mem[784] [15];
  assign _17194_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[787] [15] : \MSYNC_1r1w.synth.nz.mem[786] [15];
  assign _17195_ = \bapg_rd.w_ptr_r [1] ? _17194_ : _17193_;
  assign _17196_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[789] [15] : \MSYNC_1r1w.synth.nz.mem[788] [15];
  assign _17197_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[791] [15] : \MSYNC_1r1w.synth.nz.mem[790] [15];
  assign _17198_ = \bapg_rd.w_ptr_r [1] ? _17197_ : _17196_;
  assign _17199_ = \bapg_rd.w_ptr_r [2] ? _17198_ : _17195_;
  assign _17200_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[793] [15] : \MSYNC_1r1w.synth.nz.mem[792] [15];
  assign _17201_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[795] [15] : \MSYNC_1r1w.synth.nz.mem[794] [15];
  assign _17202_ = \bapg_rd.w_ptr_r [1] ? _17201_ : _17200_;
  assign _17203_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[797] [15] : \MSYNC_1r1w.synth.nz.mem[796] [15];
  assign _17204_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[799] [15] : \MSYNC_1r1w.synth.nz.mem[798] [15];
  assign _17205_ = \bapg_rd.w_ptr_r [1] ? _17204_ : _17203_;
  assign _17206_ = \bapg_rd.w_ptr_r [2] ? _17205_ : _17202_;
  assign _17207_ = \bapg_rd.w_ptr_r [3] ? _17206_ : _17199_;
  assign _17208_ = \bapg_rd.w_ptr_r [4] ? _17207_ : _17192_;
  assign _17209_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[801] [15] : \MSYNC_1r1w.synth.nz.mem[800] [15];
  assign _17210_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[803] [15] : \MSYNC_1r1w.synth.nz.mem[802] [15];
  assign _17211_ = \bapg_rd.w_ptr_r [1] ? _17210_ : _17209_;
  assign _17212_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[805] [15] : \MSYNC_1r1w.synth.nz.mem[804] [15];
  assign _17213_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[807] [15] : \MSYNC_1r1w.synth.nz.mem[806] [15];
  assign _17214_ = \bapg_rd.w_ptr_r [1] ? _17213_ : _17212_;
  assign _17215_ = \bapg_rd.w_ptr_r [2] ? _17214_ : _17211_;
  assign _17216_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[809] [15] : \MSYNC_1r1w.synth.nz.mem[808] [15];
  assign _17217_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[811] [15] : \MSYNC_1r1w.synth.nz.mem[810] [15];
  assign _17218_ = \bapg_rd.w_ptr_r [1] ? _17217_ : _17216_;
  assign _17219_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[813] [15] : \MSYNC_1r1w.synth.nz.mem[812] [15];
  assign _17220_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[815] [15] : \MSYNC_1r1w.synth.nz.mem[814] [15];
  assign _17221_ = \bapg_rd.w_ptr_r [1] ? _17220_ : _17219_;
  assign _17222_ = \bapg_rd.w_ptr_r [2] ? _17221_ : _17218_;
  assign _17223_ = \bapg_rd.w_ptr_r [3] ? _17222_ : _17215_;
  assign _17224_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[817] [15] : \MSYNC_1r1w.synth.nz.mem[816] [15];
  assign _17225_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[819] [15] : \MSYNC_1r1w.synth.nz.mem[818] [15];
  assign _17226_ = \bapg_rd.w_ptr_r [1] ? _17225_ : _17224_;
  assign _17227_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[821] [15] : \MSYNC_1r1w.synth.nz.mem[820] [15];
  assign _17228_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[823] [15] : \MSYNC_1r1w.synth.nz.mem[822] [15];
  assign _17229_ = \bapg_rd.w_ptr_r [1] ? _17228_ : _17227_;
  assign _17230_ = \bapg_rd.w_ptr_r [2] ? _17229_ : _17226_;
  assign _17231_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[825] [15] : \MSYNC_1r1w.synth.nz.mem[824] [15];
  assign _17232_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[827] [15] : \MSYNC_1r1w.synth.nz.mem[826] [15];
  assign _17233_ = \bapg_rd.w_ptr_r [1] ? _17232_ : _17231_;
  assign _17234_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[829] [15] : \MSYNC_1r1w.synth.nz.mem[828] [15];
  assign _17235_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[831] [15] : \MSYNC_1r1w.synth.nz.mem[830] [15];
  assign _17236_ = \bapg_rd.w_ptr_r [1] ? _17235_ : _17234_;
  assign _17237_ = \bapg_rd.w_ptr_r [2] ? _17236_ : _17233_;
  assign _17238_ = \bapg_rd.w_ptr_r [3] ? _17237_ : _17230_;
  assign _17239_ = \bapg_rd.w_ptr_r [4] ? _17238_ : _17223_;
  assign _17240_ = \bapg_rd.w_ptr_r [5] ? _17239_ : _17208_;
  assign _17241_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[833] [15] : \MSYNC_1r1w.synth.nz.mem[832] [15];
  assign _17242_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[835] [15] : \MSYNC_1r1w.synth.nz.mem[834] [15];
  assign _17243_ = \bapg_rd.w_ptr_r [1] ? _17242_ : _17241_;
  assign _17244_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[837] [15] : \MSYNC_1r1w.synth.nz.mem[836] [15];
  assign _17245_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[839] [15] : \MSYNC_1r1w.synth.nz.mem[838] [15];
  assign _17246_ = \bapg_rd.w_ptr_r [1] ? _17245_ : _17244_;
  assign _17247_ = \bapg_rd.w_ptr_r [2] ? _17246_ : _17243_;
  assign _17248_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[841] [15] : \MSYNC_1r1w.synth.nz.mem[840] [15];
  assign _17249_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[843] [15] : \MSYNC_1r1w.synth.nz.mem[842] [15];
  assign _17250_ = \bapg_rd.w_ptr_r [1] ? _17249_ : _17248_;
  assign _17251_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[845] [15] : \MSYNC_1r1w.synth.nz.mem[844] [15];
  assign _17252_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[847] [15] : \MSYNC_1r1w.synth.nz.mem[846] [15];
  assign _17253_ = \bapg_rd.w_ptr_r [1] ? _17252_ : _17251_;
  assign _17254_ = \bapg_rd.w_ptr_r [2] ? _17253_ : _17250_;
  assign _17255_ = \bapg_rd.w_ptr_r [3] ? _17254_ : _17247_;
  assign _17256_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[849] [15] : \MSYNC_1r1w.synth.nz.mem[848] [15];
  assign _17257_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[851] [15] : \MSYNC_1r1w.synth.nz.mem[850] [15];
  assign _17258_ = \bapg_rd.w_ptr_r [1] ? _17257_ : _17256_;
  assign _17259_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[853] [15] : \MSYNC_1r1w.synth.nz.mem[852] [15];
  assign _17260_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[855] [15] : \MSYNC_1r1w.synth.nz.mem[854] [15];
  assign _17261_ = \bapg_rd.w_ptr_r [1] ? _17260_ : _17259_;
  assign _17262_ = \bapg_rd.w_ptr_r [2] ? _17261_ : _17258_;
  assign _17263_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[857] [15] : \MSYNC_1r1w.synth.nz.mem[856] [15];
  assign _17264_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[859] [15] : \MSYNC_1r1w.synth.nz.mem[858] [15];
  assign _17265_ = \bapg_rd.w_ptr_r [1] ? _17264_ : _17263_;
  assign _17266_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[861] [15] : \MSYNC_1r1w.synth.nz.mem[860] [15];
  assign _17267_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[863] [15] : \MSYNC_1r1w.synth.nz.mem[862] [15];
  assign _17268_ = \bapg_rd.w_ptr_r [1] ? _17267_ : _17266_;
  assign _17269_ = \bapg_rd.w_ptr_r [2] ? _17268_ : _17265_;
  assign _17270_ = \bapg_rd.w_ptr_r [3] ? _17269_ : _17262_;
  assign _17271_ = \bapg_rd.w_ptr_r [4] ? _17270_ : _17255_;
  assign _17272_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[865] [15] : \MSYNC_1r1w.synth.nz.mem[864] [15];
  assign _17273_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[867] [15] : \MSYNC_1r1w.synth.nz.mem[866] [15];
  assign _17274_ = \bapg_rd.w_ptr_r [1] ? _17273_ : _17272_;
  assign _17275_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[869] [15] : \MSYNC_1r1w.synth.nz.mem[868] [15];
  assign _17276_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[871] [15] : \MSYNC_1r1w.synth.nz.mem[870] [15];
  assign _17277_ = \bapg_rd.w_ptr_r [1] ? _17276_ : _17275_;
  assign _17278_ = \bapg_rd.w_ptr_r [2] ? _17277_ : _17274_;
  assign _17279_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[873] [15] : \MSYNC_1r1w.synth.nz.mem[872] [15];
  assign _17280_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[875] [15] : \MSYNC_1r1w.synth.nz.mem[874] [15];
  assign _17281_ = \bapg_rd.w_ptr_r [1] ? _17280_ : _17279_;
  assign _17282_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[877] [15] : \MSYNC_1r1w.synth.nz.mem[876] [15];
  assign _17283_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[879] [15] : \MSYNC_1r1w.synth.nz.mem[878] [15];
  assign _17284_ = \bapg_rd.w_ptr_r [1] ? _17283_ : _17282_;
  assign _17285_ = \bapg_rd.w_ptr_r [2] ? _17284_ : _17281_;
  assign _17286_ = \bapg_rd.w_ptr_r [3] ? _17285_ : _17278_;
  assign _17287_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[881] [15] : \MSYNC_1r1w.synth.nz.mem[880] [15];
  assign _17288_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[883] [15] : \MSYNC_1r1w.synth.nz.mem[882] [15];
  assign _17289_ = \bapg_rd.w_ptr_r [1] ? _17288_ : _17287_;
  assign _17290_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[885] [15] : \MSYNC_1r1w.synth.nz.mem[884] [15];
  assign _17291_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[887] [15] : \MSYNC_1r1w.synth.nz.mem[886] [15];
  assign _17292_ = \bapg_rd.w_ptr_r [1] ? _17291_ : _17290_;
  assign _17293_ = \bapg_rd.w_ptr_r [2] ? _17292_ : _17289_;
  assign _17294_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[889] [15] : \MSYNC_1r1w.synth.nz.mem[888] [15];
  assign _17295_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[891] [15] : \MSYNC_1r1w.synth.nz.mem[890] [15];
  assign _17296_ = \bapg_rd.w_ptr_r [1] ? _17295_ : _17294_;
  assign _17297_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[893] [15] : \MSYNC_1r1w.synth.nz.mem[892] [15];
  assign _17298_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[895] [15] : \MSYNC_1r1w.synth.nz.mem[894] [15];
  assign _17299_ = \bapg_rd.w_ptr_r [1] ? _17298_ : _17297_;
  assign _17300_ = \bapg_rd.w_ptr_r [2] ? _17299_ : _17296_;
  assign _17301_ = \bapg_rd.w_ptr_r [3] ? _17300_ : _17293_;
  assign _17302_ = \bapg_rd.w_ptr_r [4] ? _17301_ : _17286_;
  assign _17303_ = \bapg_rd.w_ptr_r [5] ? _17302_ : _17271_;
  assign _17304_ = \bapg_rd.w_ptr_r [6] ? _17303_ : _17240_;
  assign _17305_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[897] [15] : \MSYNC_1r1w.synth.nz.mem[896] [15];
  assign _17306_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[899] [15] : \MSYNC_1r1w.synth.nz.mem[898] [15];
  assign _17307_ = \bapg_rd.w_ptr_r [1] ? _17306_ : _17305_;
  assign _17308_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[901] [15] : \MSYNC_1r1w.synth.nz.mem[900] [15];
  assign _17309_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[903] [15] : \MSYNC_1r1w.synth.nz.mem[902] [15];
  assign _17310_ = \bapg_rd.w_ptr_r [1] ? _17309_ : _17308_;
  assign _17311_ = \bapg_rd.w_ptr_r [2] ? _17310_ : _17307_;
  assign _17312_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[905] [15] : \MSYNC_1r1w.synth.nz.mem[904] [15];
  assign _17313_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[907] [15] : \MSYNC_1r1w.synth.nz.mem[906] [15];
  assign _17314_ = \bapg_rd.w_ptr_r [1] ? _17313_ : _17312_;
  assign _17315_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[909] [15] : \MSYNC_1r1w.synth.nz.mem[908] [15];
  assign _17316_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[911] [15] : \MSYNC_1r1w.synth.nz.mem[910] [15];
  assign _17317_ = \bapg_rd.w_ptr_r [1] ? _17316_ : _17315_;
  assign _17318_ = \bapg_rd.w_ptr_r [2] ? _17317_ : _17314_;
  assign _17319_ = \bapg_rd.w_ptr_r [3] ? _17318_ : _17311_;
  assign _17320_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[913] [15] : \MSYNC_1r1w.synth.nz.mem[912] [15];
  assign _17321_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[915] [15] : \MSYNC_1r1w.synth.nz.mem[914] [15];
  assign _17322_ = \bapg_rd.w_ptr_r [1] ? _17321_ : _17320_;
  assign _17323_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[917] [15] : \MSYNC_1r1w.synth.nz.mem[916] [15];
  assign _17324_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[919] [15] : \MSYNC_1r1w.synth.nz.mem[918] [15];
  assign _17325_ = \bapg_rd.w_ptr_r [1] ? _17324_ : _17323_;
  assign _17326_ = \bapg_rd.w_ptr_r [2] ? _17325_ : _17322_;
  assign _17327_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[921] [15] : \MSYNC_1r1w.synth.nz.mem[920] [15];
  assign _17328_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[923] [15] : \MSYNC_1r1w.synth.nz.mem[922] [15];
  assign _17329_ = \bapg_rd.w_ptr_r [1] ? _17328_ : _17327_;
  assign _17330_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[925] [15] : \MSYNC_1r1w.synth.nz.mem[924] [15];
  assign _17331_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[927] [15] : \MSYNC_1r1w.synth.nz.mem[926] [15];
  assign _17332_ = \bapg_rd.w_ptr_r [1] ? _17331_ : _17330_;
  assign _17333_ = \bapg_rd.w_ptr_r [2] ? _17332_ : _17329_;
  assign _17334_ = \bapg_rd.w_ptr_r [3] ? _17333_ : _17326_;
  assign _17335_ = \bapg_rd.w_ptr_r [4] ? _17334_ : _17319_;
  assign _17336_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[929] [15] : \MSYNC_1r1w.synth.nz.mem[928] [15];
  assign _17337_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[931] [15] : \MSYNC_1r1w.synth.nz.mem[930] [15];
  assign _17338_ = \bapg_rd.w_ptr_r [1] ? _17337_ : _17336_;
  assign _17339_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[933] [15] : \MSYNC_1r1w.synth.nz.mem[932] [15];
  assign _17340_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[935] [15] : \MSYNC_1r1w.synth.nz.mem[934] [15];
  assign _17341_ = \bapg_rd.w_ptr_r [1] ? _17340_ : _17339_;
  assign _17342_ = \bapg_rd.w_ptr_r [2] ? _17341_ : _17338_;
  assign _17343_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[937] [15] : \MSYNC_1r1w.synth.nz.mem[936] [15];
  assign _17344_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[939] [15] : \MSYNC_1r1w.synth.nz.mem[938] [15];
  assign _17345_ = \bapg_rd.w_ptr_r [1] ? _17344_ : _17343_;
  assign _17346_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[941] [15] : \MSYNC_1r1w.synth.nz.mem[940] [15];
  assign _17347_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[943] [15] : \MSYNC_1r1w.synth.nz.mem[942] [15];
  assign _17348_ = \bapg_rd.w_ptr_r [1] ? _17347_ : _17346_;
  assign _17349_ = \bapg_rd.w_ptr_r [2] ? _17348_ : _17345_;
  assign _17350_ = \bapg_rd.w_ptr_r [3] ? _17349_ : _17342_;
  assign _17351_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[945] [15] : \MSYNC_1r1w.synth.nz.mem[944] [15];
  assign _17352_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[947] [15] : \MSYNC_1r1w.synth.nz.mem[946] [15];
  assign _17353_ = \bapg_rd.w_ptr_r [1] ? _17352_ : _17351_;
  assign _17354_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[949] [15] : \MSYNC_1r1w.synth.nz.mem[948] [15];
  assign _17355_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[951] [15] : \MSYNC_1r1w.synth.nz.mem[950] [15];
  assign _17356_ = \bapg_rd.w_ptr_r [1] ? _17355_ : _17354_;
  assign _17357_ = \bapg_rd.w_ptr_r [2] ? _17356_ : _17353_;
  assign _17358_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[953] [15] : \MSYNC_1r1w.synth.nz.mem[952] [15];
  assign _17359_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[955] [15] : \MSYNC_1r1w.synth.nz.mem[954] [15];
  assign _17360_ = \bapg_rd.w_ptr_r [1] ? _17359_ : _17358_;
  assign _17361_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[957] [15] : \MSYNC_1r1w.synth.nz.mem[956] [15];
  assign _17362_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[959] [15] : \MSYNC_1r1w.synth.nz.mem[958] [15];
  assign _17363_ = \bapg_rd.w_ptr_r [1] ? _17362_ : _17361_;
  assign _17364_ = \bapg_rd.w_ptr_r [2] ? _17363_ : _17360_;
  assign _17365_ = \bapg_rd.w_ptr_r [3] ? _17364_ : _17357_;
  assign _17366_ = \bapg_rd.w_ptr_r [4] ? _17365_ : _17350_;
  assign _17367_ = \bapg_rd.w_ptr_r [5] ? _17366_ : _17335_;
  assign _17368_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[961] [15] : \MSYNC_1r1w.synth.nz.mem[960] [15];
  assign _17369_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[963] [15] : \MSYNC_1r1w.synth.nz.mem[962] [15];
  assign _17370_ = \bapg_rd.w_ptr_r [1] ? _17369_ : _17368_;
  assign _17371_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[965] [15] : \MSYNC_1r1w.synth.nz.mem[964] [15];
  assign _17372_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[967] [15] : \MSYNC_1r1w.synth.nz.mem[966] [15];
  assign _17373_ = \bapg_rd.w_ptr_r [1] ? _17372_ : _17371_;
  assign _17374_ = \bapg_rd.w_ptr_r [2] ? _17373_ : _17370_;
  assign _17375_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[969] [15] : \MSYNC_1r1w.synth.nz.mem[968] [15];
  assign _17376_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[971] [15] : \MSYNC_1r1w.synth.nz.mem[970] [15];
  assign _17377_ = \bapg_rd.w_ptr_r [1] ? _17376_ : _17375_;
  assign _17378_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[973] [15] : \MSYNC_1r1w.synth.nz.mem[972] [15];
  assign _17379_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[975] [15] : \MSYNC_1r1w.synth.nz.mem[974] [15];
  assign _17380_ = \bapg_rd.w_ptr_r [1] ? _17379_ : _17378_;
  assign _17381_ = \bapg_rd.w_ptr_r [2] ? _17380_ : _17377_;
  assign _17382_ = \bapg_rd.w_ptr_r [3] ? _17381_ : _17374_;
  assign _17383_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[977] [15] : \MSYNC_1r1w.synth.nz.mem[976] [15];
  assign _17384_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[979] [15] : \MSYNC_1r1w.synth.nz.mem[978] [15];
  assign _17385_ = \bapg_rd.w_ptr_r [1] ? _17384_ : _17383_;
  assign _17386_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[981] [15] : \MSYNC_1r1w.synth.nz.mem[980] [15];
  assign _17387_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[983] [15] : \MSYNC_1r1w.synth.nz.mem[982] [15];
  assign _17388_ = \bapg_rd.w_ptr_r [1] ? _17387_ : _17386_;
  assign _17389_ = \bapg_rd.w_ptr_r [2] ? _17388_ : _17385_;
  assign _17390_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[985] [15] : \MSYNC_1r1w.synth.nz.mem[984] [15];
  assign _17391_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[987] [15] : \MSYNC_1r1w.synth.nz.mem[986] [15];
  assign _17392_ = \bapg_rd.w_ptr_r [1] ? _17391_ : _17390_;
  assign _17393_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[989] [15] : \MSYNC_1r1w.synth.nz.mem[988] [15];
  assign _17394_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[991] [15] : \MSYNC_1r1w.synth.nz.mem[990] [15];
  assign _17395_ = \bapg_rd.w_ptr_r [1] ? _17394_ : _17393_;
  assign _17396_ = \bapg_rd.w_ptr_r [2] ? _17395_ : _17392_;
  assign _17397_ = \bapg_rd.w_ptr_r [3] ? _17396_ : _17389_;
  assign _17398_ = \bapg_rd.w_ptr_r [4] ? _17397_ : _17382_;
  assign _17399_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[993] [15] : \MSYNC_1r1w.synth.nz.mem[992] [15];
  assign _17400_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[995] [15] : \MSYNC_1r1w.synth.nz.mem[994] [15];
  assign _17401_ = \bapg_rd.w_ptr_r [1] ? _17400_ : _17399_;
  assign _17402_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[997] [15] : \MSYNC_1r1w.synth.nz.mem[996] [15];
  assign _17403_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[999] [15] : \MSYNC_1r1w.synth.nz.mem[998] [15];
  assign _17404_ = \bapg_rd.w_ptr_r [1] ? _17403_ : _17402_;
  assign _17405_ = \bapg_rd.w_ptr_r [2] ? _17404_ : _17401_;
  assign _17406_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1001] [15] : \MSYNC_1r1w.synth.nz.mem[1000] [15];
  assign _17407_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1003] [15] : \MSYNC_1r1w.synth.nz.mem[1002] [15];
  assign _17408_ = \bapg_rd.w_ptr_r [1] ? _17407_ : _17406_;
  assign _17409_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1005] [15] : \MSYNC_1r1w.synth.nz.mem[1004] [15];
  assign _17410_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1007] [15] : \MSYNC_1r1w.synth.nz.mem[1006] [15];
  assign _17411_ = \bapg_rd.w_ptr_r [1] ? _17410_ : _17409_;
  assign _17412_ = \bapg_rd.w_ptr_r [2] ? _17411_ : _17408_;
  assign _17413_ = \bapg_rd.w_ptr_r [3] ? _17412_ : _17405_;
  assign _17414_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1009] [15] : \MSYNC_1r1w.synth.nz.mem[1008] [15];
  assign _17415_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1011] [15] : \MSYNC_1r1w.synth.nz.mem[1010] [15];
  assign _17416_ = \bapg_rd.w_ptr_r [1] ? _17415_ : _17414_;
  assign _17417_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1013] [15] : \MSYNC_1r1w.synth.nz.mem[1012] [15];
  assign _17418_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1015] [15] : \MSYNC_1r1w.synth.nz.mem[1014] [15];
  assign _17419_ = \bapg_rd.w_ptr_r [1] ? _17418_ : _17417_;
  assign _17420_ = \bapg_rd.w_ptr_r [2] ? _17419_ : _17416_;
  assign _17421_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1017] [15] : \MSYNC_1r1w.synth.nz.mem[1016] [15];
  assign _17422_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1019] [15] : \MSYNC_1r1w.synth.nz.mem[1018] [15];
  assign _17423_ = \bapg_rd.w_ptr_r [1] ? _17422_ : _17421_;
  assign _17424_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1021] [15] : \MSYNC_1r1w.synth.nz.mem[1020] [15];
  assign _17425_ = \bapg_rd.w_ptr_r [0] ? \MSYNC_1r1w.synth.nz.mem[1023] [15] : \MSYNC_1r1w.synth.nz.mem[1022] [15];
  assign _17426_ = \bapg_rd.w_ptr_r [1] ? _17425_ : _17424_;
  assign _17427_ = \bapg_rd.w_ptr_r [2] ? _17426_ : _17423_;
  assign _17428_ = \bapg_rd.w_ptr_r [3] ? _17427_ : _17420_;
  assign _17429_ = \bapg_rd.w_ptr_r [4] ? _17428_ : _17413_;
  assign _17430_ = \bapg_rd.w_ptr_r [5] ? _17429_ : _17398_;
  assign _17431_ = \bapg_rd.w_ptr_r [6] ? _17430_ : _17367_;
  assign _17432_ = \bapg_rd.w_ptr_r [7] ? _17431_ : _17304_;
  assign _17433_ = \bapg_rd.w_ptr_r [8] ? _17432_ : _17177_;
  assign r_data_o[15] = \bapg_rd.w_ptr_r [9] ? _17433_ : _16922_;
  assign _00000_ = \bapg_wr.w_ptr_p1_r [2] ^ \bapg_wr.w_ptr_p1_r [1];
  assign _00001_ = \bapg_wr.w_ptr_p1_r [3] ^ \bapg_wr.w_ptr_p1_r [2];
  assign _00002_ = \bapg_wr.w_ptr_p1_r [4] ^ \bapg_wr.w_ptr_p1_r [3];
  assign _00003_ = \bapg_wr.w_ptr_p1_r [5] ^ \bapg_wr.w_ptr_p1_r [4];
  assign _00004_ = \bapg_wr.w_ptr_p1_r [6] ^ \bapg_wr.w_ptr_p1_r [5];
  assign _00005_ = \bapg_wr.w_ptr_p1_r [7] ^ \bapg_wr.w_ptr_p1_r [6];
  assign _00006_ = \bapg_wr.w_ptr_p1_r [8] ^ \bapg_wr.w_ptr_p1_r [7];
  assign _00007_ = \bapg_wr.w_ptr_p1_r [9] ^ \bapg_wr.w_ptr_p1_r [8];
  assign _00008_ = \bapg_wr.w_ptr_p1_r [10] ^ \bapg_wr.w_ptr_p1_r [9];
  assign _00009_ = \bapg_rd.w_ptr_p1_r [2] ^ \bapg_rd.w_ptr_p1_r [1];
  assign _00010_ = \bapg_rd.w_ptr_p1_r [3] ^ \bapg_rd.w_ptr_p1_r [2];
  assign _00011_ = \bapg_rd.w_ptr_p1_r [4] ^ \bapg_rd.w_ptr_p1_r [3];
  assign _00012_ = \bapg_rd.w_ptr_p1_r [5] ^ \bapg_rd.w_ptr_p1_r [4];
  assign _00013_ = \bapg_rd.w_ptr_p1_r [6] ^ \bapg_rd.w_ptr_p1_r [5];
  assign _00014_ = \bapg_rd.w_ptr_p1_r [7] ^ \bapg_rd.w_ptr_p1_r [6];
  assign _00015_ = \bapg_rd.w_ptr_p1_r [8] ^ \bapg_rd.w_ptr_p1_r [7];
  assign _00016_ = \bapg_rd.w_ptr_p1_r [9] ^ \bapg_rd.w_ptr_p1_r [8];
  assign _00017_ = \bapg_rd.w_ptr_p1_r [10] ^ \bapg_rd.w_ptr_p1_r [9];
  assign _17434_ = \bapg_wr.w_ptr_r [1] | \bapg_wr.w_ptr_r [0];
  assign _17435_ = \bapg_wr.w_ptr_r [4] | \bapg_wr.w_ptr_r [3];
  assign _17436_ = _17435_ | \bapg_wr.w_ptr_r [2];
  assign _17437_ = _17436_ | _17434_;
  assign _17438_ = \bapg_wr.w_ptr_r [6] | \bapg_wr.w_ptr_r [5];
  assign _17439_ = \bapg_wr.w_ptr_r [9] | \bapg_wr.w_ptr_r [8];
  assign _17440_ = _17439_ | \bapg_wr.w_ptr_r [7];
  assign _17441_ = _17440_ | _17438_;
  assign _17442_ = _17441_ | _17437_;
  assign _00018_ = w_enq_i & ~(_17442_);
  assign _17443_ = \bapg_wr.w_ptr_r [1] | ~(\bapg_wr.w_ptr_r [0]);
  assign _17444_ = _17443_ | _17436_;
  assign _17445_ = _17444_ | _17441_;
  assign _00153_ = w_enq_i & ~(_17445_);
  assign _17446_ = \bapg_wr.w_ptr_r [0] | ~(\bapg_wr.w_ptr_r [1]);
  assign _17447_ = _17446_ | _17436_;
  assign _17448_ = _17447_ | _17441_;
  assign _00264_ = w_enq_i & ~(_17448_);
  assign _17449_ = ~(\bapg_wr.w_ptr_r [1] & \bapg_wr.w_ptr_r [0]);
  assign _17450_ = _17449_ | _17436_;
  assign _17451_ = _17450_ | _17441_;
  assign _00375_ = w_enq_i & ~(_17451_);
  assign _17452_ = ~\bapg_wr.w_ptr_r [2];
  assign _17453_ = _17435_ | _17452_;
  assign _17454_ = _17453_ | _17434_;
  assign _17455_ = _17454_ | _17441_;
  assign _00486_ = w_enq_i & ~(_17455_);
  assign _17456_ = _17453_ | _17443_;
  assign _17457_ = _17456_ | _17441_;
  assign _00597_ = w_enq_i & ~(_17457_);
  assign _17458_ = _17453_ | _17446_;
  assign _17459_ = _17458_ | _17441_;
  assign _00708_ = w_enq_i & ~(_17459_);
  assign _17460_ = _17453_ | _17449_;
  assign _17461_ = _17460_ | _17441_;
  assign _00819_ = w_enq_i & ~(_17461_);
  assign _17462_ = \bapg_wr.w_ptr_r [4] | ~(\bapg_wr.w_ptr_r [3]);
  assign _17463_ = _17462_ | \bapg_wr.w_ptr_r [2];
  assign _17464_ = _17463_ | _17434_;
  assign _17465_ = _17464_ | _17441_;
  assign _00930_ = w_enq_i & ~(_17465_);
  assign _17466_ = _17463_ | _17443_;
  assign _17467_ = _17466_ | _17441_;
  assign _01041_ = w_enq_i & ~(_17467_);
  assign _17468_ = _17463_ | _17446_;
  assign _17469_ = _17468_ | _17441_;
  assign _00053_ = w_enq_i & ~(_17469_);
  assign _17470_ = _17463_ | _17449_;
  assign _17471_ = _17470_ | _17441_;
  assign _00064_ = w_enq_i & ~(_17471_);
  assign _17472_ = _17462_ | _17452_;
  assign _17473_ = _17472_ | _17434_;
  assign _17474_ = _17473_ | _17441_;
  assign _00075_ = w_enq_i & ~(_17474_);
  assign _17475_ = _17472_ | _17443_;
  assign _17476_ = _17475_ | _17441_;
  assign _00086_ = w_enq_i & ~(_17476_);
  assign _17477_ = _17472_ | _17446_;
  assign _17478_ = _17477_ | _17441_;
  assign _00097_ = w_enq_i & ~(_17478_);
  assign _17479_ = _17472_ | _17449_;
  assign _17480_ = _17479_ | _17441_;
  assign _00108_ = w_enq_i & ~(_17480_);
  assign _17481_ = \bapg_wr.w_ptr_r [3] | ~(\bapg_wr.w_ptr_r [4]);
  assign _17482_ = _17481_ | \bapg_wr.w_ptr_r [2];
  assign _17483_ = _17482_ | _17434_;
  assign _17484_ = _17483_ | _17441_;
  assign _00119_ = w_enq_i & ~(_17484_);
  assign _17485_ = _17482_ | _17443_;
  assign _17486_ = _17485_ | _17441_;
  assign _00130_ = w_enq_i & ~(_17486_);
  assign _17487_ = _17482_ | _17446_;
  assign _17488_ = _17487_ | _17441_;
  assign _00141_ = w_enq_i & ~(_17488_);
  assign _17489_ = _17482_ | _17449_;
  assign _17490_ = _17489_ | _17441_;
  assign _00152_ = w_enq_i & ~(_17490_);
  assign _17491_ = _17481_ | _17452_;
  assign _17492_ = _17491_ | _17434_;
  assign _17493_ = _17492_ | _17441_;
  assign _00164_ = w_enq_i & ~(_17493_);
  assign _17494_ = _17491_ | _17443_;
  assign _17495_ = _17494_ | _17441_;
  assign _00175_ = w_enq_i & ~(_17495_);
  assign _17496_ = _17491_ | _17446_;
  assign _17497_ = _17496_ | _17441_;
  assign _00186_ = w_enq_i & ~(_17497_);
  assign _17498_ = _17491_ | _17449_;
  assign _17499_ = _17498_ | _17441_;
  assign _00197_ = w_enq_i & ~(_17499_);
  assign _17500_ = ~(\bapg_wr.w_ptr_r [4] & \bapg_wr.w_ptr_r [3]);
  assign _17501_ = _17500_ | \bapg_wr.w_ptr_r [2];
  assign _17502_ = _17501_ | _17434_;
  assign _17503_ = _17502_ | _17441_;
  assign _00208_ = w_enq_i & ~(_17503_);
  assign _17504_ = _17501_ | _17443_;
  assign _17505_ = _17504_ | _17441_;
  assign _00219_ = w_enq_i & ~(_17505_);
  assign _17506_ = _17501_ | _17446_;
  assign _17507_ = _17506_ | _17441_;
  assign _00230_ = w_enq_i & ~(_17507_);
  assign _17508_ = _17501_ | _17449_;
  assign _17509_ = _17508_ | _17441_;
  assign _00241_ = w_enq_i & ~(_17509_);
  assign _17510_ = _17500_ | _17452_;
  assign _17511_ = _17510_ | _17434_;
  assign _17512_ = _17511_ | _17441_;
  assign _00252_ = w_enq_i & ~(_17512_);
  assign _17513_ = _17510_ | _17443_;
  assign _17514_ = _17513_ | _17441_;
  assign _00263_ = w_enq_i & ~(_17514_);
  assign _17515_ = _17510_ | _17446_;
  assign _17516_ = _17515_ | _17441_;
  assign _00275_ = w_enq_i & ~(_17516_);
  assign _17517_ = _17510_ | _17449_;
  assign _17518_ = _17517_ | _17441_;
  assign _00286_ = w_enq_i & ~(_17518_);
  assign _17519_ = \bapg_wr.w_ptr_r [6] | ~(\bapg_wr.w_ptr_r [5]);
  assign _17520_ = _17519_ | _17440_;
  assign _17521_ = _17520_ | _17437_;
  assign _00297_ = w_enq_i & ~(_17521_);
  assign _17522_ = _17520_ | _17444_;
  assign _00308_ = w_enq_i & ~(_17522_);
  assign _17523_ = _17520_ | _17447_;
  assign _00319_ = w_enq_i & ~(_17523_);
  assign _17524_ = _17520_ | _17450_;
  assign _00330_ = w_enq_i & ~(_17524_);
  assign _17525_ = _17520_ | _17454_;
  assign _00341_ = w_enq_i & ~(_17525_);
  assign _17526_ = _17520_ | _17456_;
  assign _00352_ = w_enq_i & ~(_17526_);
  assign _17527_ = _17520_ | _17458_;
  assign _00363_ = w_enq_i & ~(_17527_);
  assign _17528_ = _17520_ | _17460_;
  assign _00374_ = w_enq_i & ~(_17528_);
  assign _17529_ = _17520_ | _17464_;
  assign _00386_ = w_enq_i & ~(_17529_);
  assign _17530_ = _17520_ | _17466_;
  assign _00397_ = w_enq_i & ~(_17530_);
  assign _17531_ = _17520_ | _17468_;
  assign _00408_ = w_enq_i & ~(_17531_);
  assign _17532_ = _17520_ | _17470_;
  assign _00419_ = w_enq_i & ~(_17532_);
  assign _17533_ = _17520_ | _17473_;
  assign _00430_ = w_enq_i & ~(_17533_);
  assign _17534_ = _17520_ | _17475_;
  assign _00441_ = w_enq_i & ~(_17534_);
  assign _17535_ = _17520_ | _17477_;
  assign _00452_ = w_enq_i & ~(_17535_);
  assign _17536_ = _17520_ | _17479_;
  assign _00463_ = w_enq_i & ~(_17536_);
  assign _17537_ = _17520_ | _17483_;
  assign _00474_ = w_enq_i & ~(_17537_);
  assign _17538_ = _17520_ | _17485_;
  assign _00485_ = w_enq_i & ~(_17538_);
  assign _17539_ = _17520_ | _17487_;
  assign _00497_ = w_enq_i & ~(_17539_);
  assign _17540_ = _17520_ | _17489_;
  assign _00508_ = w_enq_i & ~(_17540_);
  assign _17541_ = _17520_ | _17492_;
  assign _00519_ = w_enq_i & ~(_17541_);
  assign _17542_ = _17520_ | _17494_;
  assign _00530_ = w_enq_i & ~(_17542_);
  assign _17543_ = _17520_ | _17496_;
  assign _00541_ = w_enq_i & ~(_17543_);
  assign _17544_ = _17520_ | _17498_;
  assign _00552_ = w_enq_i & ~(_17544_);
  assign _17545_ = _17520_ | _17502_;
  assign _00563_ = w_enq_i & ~(_17545_);
  assign _17546_ = _17520_ | _17504_;
  assign _00574_ = w_enq_i & ~(_17546_);
  assign _17547_ = _17520_ | _17506_;
  assign _00585_ = w_enq_i & ~(_17547_);
  assign _17548_ = _17520_ | _17508_;
  assign _00596_ = w_enq_i & ~(_17548_);
  assign _17549_ = _17520_ | _17511_;
  assign _00608_ = w_enq_i & ~(_17549_);
  assign _17550_ = _17520_ | _17513_;
  assign _00619_ = w_enq_i & ~(_17550_);
  assign _17551_ = _17520_ | _17515_;
  assign _00630_ = w_enq_i & ~(_17551_);
  assign _17552_ = _17520_ | _17517_;
  assign _00641_ = w_enq_i & ~(_17552_);
  assign _17553_ = \bapg_wr.w_ptr_r [5] | ~(\bapg_wr.w_ptr_r [6]);
  assign _17554_ = _17553_ | _17440_;
  assign _17555_ = _17554_ | _17437_;
  assign _00652_ = w_enq_i & ~(_17555_);
  assign _17556_ = _17554_ | _17444_;
  assign _00663_ = w_enq_i & ~(_17556_);
  assign _17557_ = _17554_ | _17447_;
  assign _00674_ = w_enq_i & ~(_17557_);
  assign _17558_ = _17554_ | _17450_;
  assign _00685_ = w_enq_i & ~(_17558_);
  assign _17559_ = _17554_ | _17454_;
  assign _00696_ = w_enq_i & ~(_17559_);
  assign _17560_ = _17554_ | _17456_;
  assign _00707_ = w_enq_i & ~(_17560_);
  assign _17561_ = _17554_ | _17458_;
  assign _00719_ = w_enq_i & ~(_17561_);
  assign _17562_ = _17554_ | _17460_;
  assign _00730_ = w_enq_i & ~(_17562_);
  assign _17563_ = _17554_ | _17464_;
  assign _00741_ = w_enq_i & ~(_17563_);
  assign _17564_ = _17554_ | _17466_;
  assign _00752_ = w_enq_i & ~(_17564_);
  assign _17565_ = _17554_ | _17468_;
  assign _00763_ = w_enq_i & ~(_17565_);
  assign _17566_ = _17554_ | _17470_;
  assign _00774_ = w_enq_i & ~(_17566_);
  assign _17567_ = _17554_ | _17473_;
  assign _00785_ = w_enq_i & ~(_17567_);
  assign _17568_ = _17554_ | _17475_;
  assign _00796_ = w_enq_i & ~(_17568_);
  assign _17569_ = _17554_ | _17477_;
  assign _00807_ = w_enq_i & ~(_17569_);
  assign _17570_ = _17554_ | _17479_;
  assign _00818_ = w_enq_i & ~(_17570_);
  assign _17571_ = _17554_ | _17483_;
  assign _00830_ = w_enq_i & ~(_17571_);
  assign _17572_ = _17554_ | _17485_;
  assign _00841_ = w_enq_i & ~(_17572_);
  assign _17573_ = _17554_ | _17487_;
  assign _00852_ = w_enq_i & ~(_17573_);
  assign _17574_ = _17554_ | _17489_;
  assign _00863_ = w_enq_i & ~(_17574_);
  assign _17575_ = _17554_ | _17492_;
  assign _00874_ = w_enq_i & ~(_17575_);
  assign _17576_ = _17554_ | _17494_;
  assign _00885_ = w_enq_i & ~(_17576_);
  assign _17577_ = _17554_ | _17496_;
  assign _00896_ = w_enq_i & ~(_17577_);
  assign _17578_ = _17554_ | _17498_;
  assign _00907_ = w_enq_i & ~(_17578_);
  assign _17579_ = _17554_ | _17502_;
  assign _00918_ = w_enq_i & ~(_17579_);
  assign _17580_ = _17554_ | _17504_;
  assign _00929_ = w_enq_i & ~(_17580_);
  assign _17581_ = _17554_ | _17506_;
  assign _00941_ = w_enq_i & ~(_17581_);
  assign _17582_ = _17554_ | _17508_;
  assign _00952_ = w_enq_i & ~(_17582_);
  assign _17583_ = _17554_ | _17511_;
  assign _00963_ = w_enq_i & ~(_17583_);
  assign _17584_ = _17554_ | _17513_;
  assign _00974_ = w_enq_i & ~(_17584_);
  assign _17585_ = _17554_ | _17515_;
  assign _00985_ = w_enq_i & ~(_17585_);
  assign _17586_ = _17554_ | _17517_;
  assign _00996_ = w_enq_i & ~(_17586_);
  assign _17587_ = ~(\bapg_wr.w_ptr_r [6] & \bapg_wr.w_ptr_r [5]);
  assign _17588_ = _17587_ | _17440_;
  assign _17589_ = _17588_ | _17437_;
  assign _01007_ = w_enq_i & ~(_17589_);
  assign _17590_ = _17588_ | _17444_;
  assign _01018_ = w_enq_i & ~(_17590_);
  assign _17591_ = _17588_ | _17447_;
  assign _01029_ = w_enq_i & ~(_17591_);
  assign _17592_ = _17588_ | _17450_;
  assign _01040_ = w_enq_i & ~(_17592_);
  assign _17593_ = _17588_ | _17454_;
  assign _00029_ = w_enq_i & ~(_17593_);
  assign _17594_ = _17588_ | _17456_;
  assign _00040_ = w_enq_i & ~(_17594_);
  assign _17595_ = _17588_ | _17458_;
  assign _00045_ = w_enq_i & ~(_17595_);
  assign _17596_ = _17588_ | _17460_;
  assign _00046_ = w_enq_i & ~(_17596_);
  assign _17597_ = _17588_ | _17464_;
  assign _00047_ = w_enq_i & ~(_17597_);
  assign _17598_ = _17588_ | _17466_;
  assign _00048_ = w_enq_i & ~(_17598_);
  assign _17599_ = _17588_ | _17468_;
  assign _00049_ = w_enq_i & ~(_17599_);
  assign _17600_ = _17588_ | _17470_;
  assign _00050_ = w_enq_i & ~(_17600_);
  assign _17601_ = _17588_ | _17473_;
  assign _00051_ = w_enq_i & ~(_17601_);
  assign _17602_ = _17588_ | _17475_;
  assign _00052_ = w_enq_i & ~(_17602_);
  assign _17603_ = _17588_ | _17477_;
  assign _00054_ = w_enq_i & ~(_17603_);
  assign _17604_ = _17588_ | _17479_;
  assign _00055_ = w_enq_i & ~(_17604_);
  assign _17605_ = _17588_ | _17483_;
  assign _00056_ = w_enq_i & ~(_17605_);
  assign _17606_ = _17588_ | _17485_;
  assign _00057_ = w_enq_i & ~(_17606_);
  assign _17607_ = _17588_ | _17487_;
  assign _00058_ = w_enq_i & ~(_17607_);
  assign _17608_ = _17588_ | _17489_;
  assign _00059_ = w_enq_i & ~(_17608_);
  assign _17609_ = _17588_ | _17492_;
  assign _00060_ = w_enq_i & ~(_17609_);
  assign _17610_ = _17588_ | _17494_;
  assign _00061_ = w_enq_i & ~(_17610_);
  assign _17611_ = _17588_ | _17496_;
  assign _00062_ = w_enq_i & ~(_17611_);
  assign _17612_ = _17588_ | _17498_;
  assign _00063_ = w_enq_i & ~(_17612_);
  assign _17613_ = _17588_ | _17502_;
  assign _00065_ = w_enq_i & ~(_17613_);
  assign _17614_ = _17588_ | _17504_;
  assign _00066_ = w_enq_i & ~(_17614_);
  assign _17615_ = _17588_ | _17506_;
  assign _00067_ = w_enq_i & ~(_17615_);
  assign _17616_ = _17588_ | _17508_;
  assign _00068_ = w_enq_i & ~(_17616_);
  assign _17617_ = _17588_ | _17511_;
  assign _00069_ = w_enq_i & ~(_17617_);
  assign _17618_ = _17588_ | _17513_;
  assign _00070_ = w_enq_i & ~(_17618_);
  assign _17619_ = _17588_ | _17515_;
  assign _00071_ = w_enq_i & ~(_17619_);
  assign _17620_ = _17588_ | _17517_;
  assign _00072_ = w_enq_i & ~(_17620_);
  assign _17621_ = ~\bapg_wr.w_ptr_r [7];
  assign _17622_ = _17439_ | _17621_;
  assign _17623_ = _17622_ | _17438_;
  assign _17624_ = _17623_ | _17437_;
  assign _00073_ = w_enq_i & ~(_17624_);
  assign _17625_ = _17623_ | _17444_;
  assign _00074_ = w_enq_i & ~(_17625_);
  assign _17626_ = _17623_ | _17447_;
  assign _00076_ = w_enq_i & ~(_17626_);
  assign _17627_ = _17623_ | _17450_;
  assign _00077_ = w_enq_i & ~(_17627_);
  assign _17628_ = _17623_ | _17454_;
  assign _00078_ = w_enq_i & ~(_17628_);
  assign _17629_ = _17623_ | _17456_;
  assign _00079_ = w_enq_i & ~(_17629_);
  assign _17630_ = _17623_ | _17458_;
  assign _00080_ = w_enq_i & ~(_17630_);
  assign _17631_ = _17623_ | _17460_;
  assign _00081_ = w_enq_i & ~(_17631_);
  assign _17632_ = _17623_ | _17464_;
  assign _00082_ = w_enq_i & ~(_17632_);
  assign _17633_ = _17623_ | _17466_;
  assign _00083_ = w_enq_i & ~(_17633_);
  assign _17634_ = _17623_ | _17468_;
  assign _00084_ = w_enq_i & ~(_17634_);
  assign _17635_ = _17623_ | _17470_;
  assign _00085_ = w_enq_i & ~(_17635_);
  assign _17636_ = _17623_ | _17473_;
  assign _00087_ = w_enq_i & ~(_17636_);
  assign _17637_ = _17623_ | _17475_;
  assign _00088_ = w_enq_i & ~(_17637_);
  assign _17638_ = _17623_ | _17477_;
  assign _00089_ = w_enq_i & ~(_17638_);
  assign _17639_ = _17623_ | _17479_;
  assign _00090_ = w_enq_i & ~(_17639_);
  assign _17640_ = _17623_ | _17483_;
  assign _00091_ = w_enq_i & ~(_17640_);
  assign _17641_ = _17623_ | _17485_;
  assign _00092_ = w_enq_i & ~(_17641_);
  assign _17642_ = _17623_ | _17487_;
  assign _00093_ = w_enq_i & ~(_17642_);
  assign _17643_ = _17623_ | _17489_;
  assign _00094_ = w_enq_i & ~(_17643_);
  assign _17644_ = _17623_ | _17492_;
  assign _00095_ = w_enq_i & ~(_17644_);
  assign _17645_ = _17623_ | _17494_;
  assign _00096_ = w_enq_i & ~(_17645_);
  assign _17646_ = _17623_ | _17496_;
  assign _00098_ = w_enq_i & ~(_17646_);
  assign _17647_ = _17623_ | _17498_;
  assign _00099_ = w_enq_i & ~(_17647_);
  assign _17648_ = _17623_ | _17502_;
  assign _00100_ = w_enq_i & ~(_17648_);
  assign _17649_ = _17623_ | _17504_;
  assign _00101_ = w_enq_i & ~(_17649_);
  assign _17650_ = _17623_ | _17506_;
  assign _00102_ = w_enq_i & ~(_17650_);
  assign _17651_ = _17623_ | _17508_;
  assign _00103_ = w_enq_i & ~(_17651_);
  assign _17652_ = _17623_ | _17511_;
  assign _00104_ = w_enq_i & ~(_17652_);
  assign _17653_ = _17623_ | _17513_;
  assign _00105_ = w_enq_i & ~(_17653_);
  assign _17654_ = _17623_ | _17515_;
  assign _00106_ = w_enq_i & ~(_17654_);
  assign _17655_ = _17623_ | _17517_;
  assign _00107_ = w_enq_i & ~(_17655_);
  assign _17656_ = _17622_ | _17519_;
  assign _17657_ = _17656_ | _17437_;
  assign _00109_ = w_enq_i & ~(_17657_);
  assign _17658_ = _17656_ | _17444_;
  assign _00110_ = w_enq_i & ~(_17658_);
  assign _17659_ = _17656_ | _17447_;
  assign _00111_ = w_enq_i & ~(_17659_);
  assign _17660_ = _17656_ | _17450_;
  assign _00112_ = w_enq_i & ~(_17660_);
  assign _17661_ = _17656_ | _17454_;
  assign _00113_ = w_enq_i & ~(_17661_);
  assign _17662_ = _17656_ | _17456_;
  assign _00114_ = w_enq_i & ~(_17662_);
  assign _17663_ = _17656_ | _17458_;
  assign _00115_ = w_enq_i & ~(_17663_);
  assign _17664_ = _17656_ | _17460_;
  assign _00116_ = w_enq_i & ~(_17664_);
  assign _17665_ = _17656_ | _17464_;
  assign _00117_ = w_enq_i & ~(_17665_);
  assign _17666_ = _17656_ | _17466_;
  assign _00118_ = w_enq_i & ~(_17666_);
  assign _17667_ = _17656_ | _17468_;
  assign _00120_ = w_enq_i & ~(_17667_);
  assign _17668_ = _17656_ | _17470_;
  assign _00121_ = w_enq_i & ~(_17668_);
  assign _17669_ = _17656_ | _17473_;
  assign _00122_ = w_enq_i & ~(_17669_);
  assign _17670_ = _17656_ | _17475_;
  assign _00123_ = w_enq_i & ~(_17670_);
  assign _17671_ = _17656_ | _17477_;
  assign _00124_ = w_enq_i & ~(_17671_);
  assign _17672_ = _17656_ | _17479_;
  assign _00125_ = w_enq_i & ~(_17672_);
  assign _17673_ = _17656_ | _17483_;
  assign _00126_ = w_enq_i & ~(_17673_);
  assign _17674_ = _17656_ | _17485_;
  assign _00127_ = w_enq_i & ~(_17674_);
  assign _17675_ = _17656_ | _17487_;
  assign _00128_ = w_enq_i & ~(_17675_);
  assign _17676_ = _17656_ | _17489_;
  assign _00129_ = w_enq_i & ~(_17676_);
  assign _17677_ = _17656_ | _17492_;
  assign _00131_ = w_enq_i & ~(_17677_);
  assign _17678_ = _17656_ | _17494_;
  assign _00132_ = w_enq_i & ~(_17678_);
  assign _17679_ = _17656_ | _17496_;
  assign _00133_ = w_enq_i & ~(_17679_);
  assign _17680_ = _17656_ | _17498_;
  assign _00134_ = w_enq_i & ~(_17680_);
  assign _17681_ = _17656_ | _17502_;
  assign _00135_ = w_enq_i & ~(_17681_);
  assign _17682_ = _17656_ | _17504_;
  assign _00136_ = w_enq_i & ~(_17682_);
  assign _17683_ = _17656_ | _17506_;
  assign _00137_ = w_enq_i & ~(_17683_);
  assign _17684_ = _17656_ | _17508_;
  assign _00138_ = w_enq_i & ~(_17684_);
  assign _17685_ = _17656_ | _17511_;
  assign _00139_ = w_enq_i & ~(_17685_);
  assign _17686_ = _17656_ | _17513_;
  assign _00140_ = w_enq_i & ~(_17686_);
  assign _17687_ = _17656_ | _17515_;
  assign _00142_ = w_enq_i & ~(_17687_);
  assign _17688_ = _17656_ | _17517_;
  assign _00143_ = w_enq_i & ~(_17688_);
  assign _17689_ = _17622_ | _17553_;
  assign _17690_ = _17689_ | _17437_;
  assign _00144_ = w_enq_i & ~(_17690_);
  assign _17691_ = _17689_ | _17444_;
  assign _00145_ = w_enq_i & ~(_17691_);
  assign _17692_ = _17689_ | _17447_;
  assign _00146_ = w_enq_i & ~(_17692_);
  assign _17693_ = _17689_ | _17450_;
  assign _00147_ = w_enq_i & ~(_17693_);
  assign _17694_ = _17689_ | _17454_;
  assign _00148_ = w_enq_i & ~(_17694_);
  assign _17695_ = _17689_ | _17456_;
  assign _00149_ = w_enq_i & ~(_17695_);
  assign _17696_ = _17689_ | _17458_;
  assign _00150_ = w_enq_i & ~(_17696_);
  assign _17697_ = _17689_ | _17460_;
  assign _00151_ = w_enq_i & ~(_17697_);
  assign _17698_ = _17689_ | _17464_;
  assign _00154_ = w_enq_i & ~(_17698_);
  assign _17699_ = _17689_ | _17466_;
  assign _00155_ = w_enq_i & ~(_17699_);
  assign _17700_ = _17689_ | _17468_;
  assign _00156_ = w_enq_i & ~(_17700_);
  assign _17701_ = _17689_ | _17470_;
  assign _00157_ = w_enq_i & ~(_17701_);
  assign _17702_ = _17689_ | _17473_;
  assign _00158_ = w_enq_i & ~(_17702_);
  assign _17703_ = _17689_ | _17475_;
  assign _00159_ = w_enq_i & ~(_17703_);
  assign _17704_ = _17689_ | _17477_;
  assign _00160_ = w_enq_i & ~(_17704_);
  assign _17705_ = _17689_ | _17479_;
  assign _00161_ = w_enq_i & ~(_17705_);
  assign _17706_ = _17689_ | _17483_;
  assign _00162_ = w_enq_i & ~(_17706_);
  assign _17707_ = _17689_ | _17485_;
  assign _00163_ = w_enq_i & ~(_17707_);
  assign _17708_ = _17689_ | _17487_;
  assign _00165_ = w_enq_i & ~(_17708_);
  assign _17709_ = _17689_ | _17489_;
  assign _00166_ = w_enq_i & ~(_17709_);
  assign _17710_ = _17689_ | _17492_;
  assign _00167_ = w_enq_i & ~(_17710_);
  assign _17711_ = _17689_ | _17494_;
  assign _00168_ = w_enq_i & ~(_17711_);
  assign _17712_ = _17689_ | _17496_;
  assign _00169_ = w_enq_i & ~(_17712_);
  assign _17713_ = _17689_ | _17498_;
  assign _00170_ = w_enq_i & ~(_17713_);
  assign _17714_ = _17689_ | _17502_;
  assign _00171_ = w_enq_i & ~(_17714_);
  assign _17715_ = _17689_ | _17504_;
  assign _00172_ = w_enq_i & ~(_17715_);
  assign _17716_ = _17689_ | _17506_;
  assign _00173_ = w_enq_i & ~(_17716_);
  assign _17717_ = _17689_ | _17508_;
  assign _00174_ = w_enq_i & ~(_17717_);
  assign _17718_ = _17689_ | _17511_;
  assign _00176_ = w_enq_i & ~(_17718_);
  assign _17719_ = _17689_ | _17513_;
  assign _00177_ = w_enq_i & ~(_17719_);
  assign _17720_ = _17689_ | _17515_;
  assign _00178_ = w_enq_i & ~(_17720_);
  assign _17721_ = _17689_ | _17517_;
  assign _00179_ = w_enq_i & ~(_17721_);
  assign _17722_ = _17622_ | _17587_;
  assign _17723_ = _17722_ | _17437_;
  assign _00180_ = w_enq_i & ~(_17723_);
  assign _17724_ = _17722_ | _17444_;
  assign _00181_ = w_enq_i & ~(_17724_);
  assign _17725_ = _17722_ | _17447_;
  assign _00182_ = w_enq_i & ~(_17725_);
  assign _17726_ = _17722_ | _17450_;
  assign _00183_ = w_enq_i & ~(_17726_);
  assign _17727_ = _17722_ | _17454_;
  assign _00184_ = w_enq_i & ~(_17727_);
  assign _17728_ = _17722_ | _17456_;
  assign _00185_ = w_enq_i & ~(_17728_);
  assign _17729_ = _17722_ | _17458_;
  assign _00187_ = w_enq_i & ~(_17729_);
  assign _17730_ = _17722_ | _17460_;
  assign _00188_ = w_enq_i & ~(_17730_);
  assign _17731_ = _17722_ | _17464_;
  assign _00189_ = w_enq_i & ~(_17731_);
  assign _17732_ = _17722_ | _17466_;
  assign _00190_ = w_enq_i & ~(_17732_);
  assign _17733_ = _17722_ | _17468_;
  assign _00191_ = w_enq_i & ~(_17733_);
  assign _17734_ = _17722_ | _17470_;
  assign _00192_ = w_enq_i & ~(_17734_);
  assign _17735_ = _17722_ | _17473_;
  assign _00193_ = w_enq_i & ~(_17735_);
  assign _17736_ = _17722_ | _17475_;
  assign _00194_ = w_enq_i & ~(_17736_);
  assign _17737_ = _17722_ | _17477_;
  assign _00195_ = w_enq_i & ~(_17737_);
  assign _17738_ = _17722_ | _17479_;
  assign _00196_ = w_enq_i & ~(_17738_);
  assign _17739_ = _17722_ | _17483_;
  assign _00198_ = w_enq_i & ~(_17739_);
  assign _17740_ = _17722_ | _17485_;
  assign _00199_ = w_enq_i & ~(_17740_);
  assign _17741_ = _17722_ | _17487_;
  assign _00200_ = w_enq_i & ~(_17741_);
  assign _17742_ = _17722_ | _17489_;
  assign _00201_ = w_enq_i & ~(_17742_);
  assign _17743_ = _17722_ | _17492_;
  assign _00202_ = w_enq_i & ~(_17743_);
  assign _17744_ = _17722_ | _17494_;
  assign _00203_ = w_enq_i & ~(_17744_);
  assign _17745_ = _17722_ | _17496_;
  assign _00204_ = w_enq_i & ~(_17745_);
  assign _17746_ = _17722_ | _17498_;
  assign _00205_ = w_enq_i & ~(_17746_);
  assign _17747_ = _17722_ | _17502_;
  assign _00206_ = w_enq_i & ~(_17747_);
  assign _17748_ = _17722_ | _17504_;
  assign _00207_ = w_enq_i & ~(_17748_);
  assign _17749_ = _17722_ | _17506_;
  assign _00209_ = w_enq_i & ~(_17749_);
  assign _17750_ = _17722_ | _17508_;
  assign _00210_ = w_enq_i & ~(_17750_);
  assign _17751_ = _17722_ | _17511_;
  assign _00211_ = w_enq_i & ~(_17751_);
  assign _17752_ = _17722_ | _17513_;
  assign _00212_ = w_enq_i & ~(_17752_);
  assign _17753_ = _17722_ | _17515_;
  assign _00213_ = w_enq_i & ~(_17753_);
  assign _17754_ = _17722_ | _17517_;
  assign _00214_ = w_enq_i & ~(_17754_);
  assign _17755_ = \bapg_wr.w_ptr_r [9] | ~(\bapg_wr.w_ptr_r [8]);
  assign _17756_ = _17755_ | \bapg_wr.w_ptr_r [7];
  assign _17757_ = _17756_ | _17438_;
  assign _17758_ = _17757_ | _17437_;
  assign _00215_ = w_enq_i & ~(_17758_);
  assign _17759_ = _17757_ | _17444_;
  assign _00216_ = w_enq_i & ~(_17759_);
  assign _17760_ = _17757_ | _17447_;
  assign _00217_ = w_enq_i & ~(_17760_);
  assign _17761_ = _17757_ | _17450_;
  assign _00218_ = w_enq_i & ~(_17761_);
  assign _17762_ = _17757_ | _17454_;
  assign _00220_ = w_enq_i & ~(_17762_);
  assign _17763_ = _17757_ | _17456_;
  assign _00221_ = w_enq_i & ~(_17763_);
  assign _17764_ = _17757_ | _17458_;
  assign _00222_ = w_enq_i & ~(_17764_);
  assign _17765_ = _17757_ | _17460_;
  assign _00223_ = w_enq_i & ~(_17765_);
  assign _17766_ = _17757_ | _17464_;
  assign _00224_ = w_enq_i & ~(_17766_);
  assign _17767_ = _17757_ | _17466_;
  assign _00225_ = w_enq_i & ~(_17767_);
  assign _17768_ = _17757_ | _17468_;
  assign _00226_ = w_enq_i & ~(_17768_);
  assign _17769_ = _17757_ | _17470_;
  assign _00227_ = w_enq_i & ~(_17769_);
  assign _17770_ = _17757_ | _17473_;
  assign _00228_ = w_enq_i & ~(_17770_);
  assign _17771_ = _17757_ | _17475_;
  assign _00229_ = w_enq_i & ~(_17771_);
  assign _17772_ = _17757_ | _17477_;
  assign _00231_ = w_enq_i & ~(_17772_);
  assign _17773_ = _17757_ | _17479_;
  assign _00232_ = w_enq_i & ~(_17773_);
  assign _17774_ = _17757_ | _17483_;
  assign _00233_ = w_enq_i & ~(_17774_);
  assign _17775_ = _17757_ | _17485_;
  assign _00234_ = w_enq_i & ~(_17775_);
  assign _17776_ = _17757_ | _17487_;
  assign _00235_ = w_enq_i & ~(_17776_);
  assign _17777_ = _17757_ | _17489_;
  assign _00236_ = w_enq_i & ~(_17777_);
  assign _17778_ = _17757_ | _17492_;
  assign _00237_ = w_enq_i & ~(_17778_);
  assign _17779_ = _17757_ | _17494_;
  assign _00238_ = w_enq_i & ~(_17779_);
  assign _17780_ = _17757_ | _17496_;
  assign _00239_ = w_enq_i & ~(_17780_);
  assign _17781_ = _17757_ | _17498_;
  assign _00240_ = w_enq_i & ~(_17781_);
  assign _17782_ = _17757_ | _17502_;
  assign _00242_ = w_enq_i & ~(_17782_);
  assign _17783_ = _17757_ | _17504_;
  assign _00243_ = w_enq_i & ~(_17783_);
  assign _17784_ = _17757_ | _17506_;
  assign _00244_ = w_enq_i & ~(_17784_);
  assign _17785_ = _17757_ | _17508_;
  assign _00245_ = w_enq_i & ~(_17785_);
  assign _17786_ = _17757_ | _17511_;
  assign _00246_ = w_enq_i & ~(_17786_);
  assign _17787_ = _17757_ | _17513_;
  assign _00247_ = w_enq_i & ~(_17787_);
  assign _17788_ = _17757_ | _17515_;
  assign _00248_ = w_enq_i & ~(_17788_);
  assign _17789_ = _17757_ | _17517_;
  assign _00249_ = w_enq_i & ~(_17789_);
  assign _17790_ = _17756_ | _17519_;
  assign _17791_ = _17790_ | _17437_;
  assign _00250_ = w_enq_i & ~(_17791_);
  assign _17792_ = _17790_ | _17444_;
  assign _00251_ = w_enq_i & ~(_17792_);
  assign _17793_ = _17790_ | _17447_;
  assign _00253_ = w_enq_i & ~(_17793_);
  assign _17794_ = _17790_ | _17450_;
  assign _00254_ = w_enq_i & ~(_17794_);
  assign _17795_ = _17790_ | _17454_;
  assign _00255_ = w_enq_i & ~(_17795_);
  assign _17796_ = _17790_ | _17456_;
  assign _00256_ = w_enq_i & ~(_17796_);
  assign _17797_ = _17790_ | _17458_;
  assign _00257_ = w_enq_i & ~(_17797_);
  assign _17798_ = _17790_ | _17460_;
  assign _00258_ = w_enq_i & ~(_17798_);
  assign _17799_ = _17790_ | _17464_;
  assign _00259_ = w_enq_i & ~(_17799_);
  assign _17800_ = _17790_ | _17466_;
  assign _00260_ = w_enq_i & ~(_17800_);
  assign _17801_ = _17790_ | _17468_;
  assign _00261_ = w_enq_i & ~(_17801_);
  assign _17802_ = _17790_ | _17470_;
  assign _00262_ = w_enq_i & ~(_17802_);
  assign _17803_ = _17790_ | _17473_;
  assign _00265_ = w_enq_i & ~(_17803_);
  assign _17804_ = _17790_ | _17475_;
  assign _00266_ = w_enq_i & ~(_17804_);
  assign _17805_ = _17790_ | _17477_;
  assign _00267_ = w_enq_i & ~(_17805_);
  assign _17806_ = _17790_ | _17479_;
  assign _00268_ = w_enq_i & ~(_17806_);
  assign _17807_ = _17790_ | _17483_;
  assign _00269_ = w_enq_i & ~(_17807_);
  assign _17808_ = _17790_ | _17485_;
  assign _00270_ = w_enq_i & ~(_17808_);
  assign _17809_ = _17790_ | _17487_;
  assign _00271_ = w_enq_i & ~(_17809_);
  assign _17810_ = _17790_ | _17489_;
  assign _00272_ = w_enq_i & ~(_17810_);
  assign _17811_ = _17790_ | _17492_;
  assign _00273_ = w_enq_i & ~(_17811_);
  assign _17812_ = _17790_ | _17494_;
  assign _00274_ = w_enq_i & ~(_17812_);
  assign _17813_ = _17790_ | _17496_;
  assign _00276_ = w_enq_i & ~(_17813_);
  assign _17814_ = _17790_ | _17498_;
  assign _00277_ = w_enq_i & ~(_17814_);
  assign _17815_ = _17790_ | _17502_;
  assign _00278_ = w_enq_i & ~(_17815_);
  assign _17816_ = _17790_ | _17504_;
  assign _00279_ = w_enq_i & ~(_17816_);
  assign _17817_ = _17790_ | _17506_;
  assign _00280_ = w_enq_i & ~(_17817_);
  assign _17818_ = _17790_ | _17508_;
  assign _00281_ = w_enq_i & ~(_17818_);
  assign _17819_ = _17790_ | _17511_;
  assign _00282_ = w_enq_i & ~(_17819_);
  assign _17820_ = _17790_ | _17513_;
  assign _00283_ = w_enq_i & ~(_17820_);
  assign _17821_ = _17790_ | _17515_;
  assign _00284_ = w_enq_i & ~(_17821_);
  assign _17822_ = _17790_ | _17517_;
  assign _00285_ = w_enq_i & ~(_17822_);
  assign _17823_ = _17756_ | _17553_;
  assign _17824_ = _17823_ | _17437_;
  assign _00287_ = w_enq_i & ~(_17824_);
  assign _17825_ = _17823_ | _17444_;
  assign _00288_ = w_enq_i & ~(_17825_);
  assign _17826_ = _17823_ | _17447_;
  assign _00289_ = w_enq_i & ~(_17826_);
  assign _17827_ = _17823_ | _17450_;
  assign _00290_ = w_enq_i & ~(_17827_);
  assign _17828_ = _17823_ | _17454_;
  assign _00291_ = w_enq_i & ~(_17828_);
  assign _17829_ = _17823_ | _17456_;
  assign _00292_ = w_enq_i & ~(_17829_);
  assign _17830_ = _17823_ | _17458_;
  assign _00293_ = w_enq_i & ~(_17830_);
  assign _17831_ = _17823_ | _17460_;
  assign _00294_ = w_enq_i & ~(_17831_);
  assign _17832_ = _17823_ | _17464_;
  assign _00295_ = w_enq_i & ~(_17832_);
  assign _17833_ = _17823_ | _17466_;
  assign _00296_ = w_enq_i & ~(_17833_);
  assign _17834_ = _17823_ | _17468_;
  assign _00298_ = w_enq_i & ~(_17834_);
  assign _17835_ = _17823_ | _17470_;
  assign _00299_ = w_enq_i & ~(_17835_);
  assign _17836_ = _17823_ | _17473_;
  assign _00300_ = w_enq_i & ~(_17836_);
  assign _17837_ = _17823_ | _17475_;
  assign _00301_ = w_enq_i & ~(_17837_);
  assign _17838_ = _17823_ | _17477_;
  assign _00302_ = w_enq_i & ~(_17838_);
  assign _17839_ = _17823_ | _17479_;
  assign _00303_ = w_enq_i & ~(_17839_);
  assign _17840_ = _17823_ | _17483_;
  assign _00304_ = w_enq_i & ~(_17840_);
  assign _17841_ = _17823_ | _17485_;
  assign _00305_ = w_enq_i & ~(_17841_);
  assign _17842_ = _17823_ | _17487_;
  assign _00306_ = w_enq_i & ~(_17842_);
  assign _17843_ = _17823_ | _17489_;
  assign _00307_ = w_enq_i & ~(_17843_);
  assign _17844_ = _17823_ | _17492_;
  assign _00309_ = w_enq_i & ~(_17844_);
  assign _17845_ = _17823_ | _17494_;
  assign _00310_ = w_enq_i & ~(_17845_);
  assign _17846_ = _17823_ | _17496_;
  assign _00311_ = w_enq_i & ~(_17846_);
  assign _17847_ = _17823_ | _17498_;
  assign _00312_ = w_enq_i & ~(_17847_);
  assign _17848_ = _17823_ | _17502_;
  assign _00313_ = w_enq_i & ~(_17848_);
  assign _17849_ = _17823_ | _17504_;
  assign _00314_ = w_enq_i & ~(_17849_);
  assign _17850_ = _17823_ | _17506_;
  assign _00315_ = w_enq_i & ~(_17850_);
  assign _17851_ = _17823_ | _17508_;
  assign _00316_ = w_enq_i & ~(_17851_);
  assign _17852_ = _17823_ | _17511_;
  assign _00317_ = w_enq_i & ~(_17852_);
  assign _17853_ = _17823_ | _17513_;
  assign _00318_ = w_enq_i & ~(_17853_);
  assign _17854_ = _17823_ | _17515_;
  assign _00320_ = w_enq_i & ~(_17854_);
  assign _17855_ = _17823_ | _17517_;
  assign _00321_ = w_enq_i & ~(_17855_);
  assign _17856_ = _17756_ | _17587_;
  assign _17857_ = _17856_ | _17437_;
  assign _00322_ = w_enq_i & ~(_17857_);
  assign _17858_ = _17856_ | _17444_;
  assign _00323_ = w_enq_i & ~(_17858_);
  assign _17859_ = _17856_ | _17447_;
  assign _00324_ = w_enq_i & ~(_17859_);
  assign _17860_ = _17856_ | _17450_;
  assign _00325_ = w_enq_i & ~(_17860_);
  assign _17861_ = _17856_ | _17454_;
  assign _00326_ = w_enq_i & ~(_17861_);
  assign _17862_ = _17856_ | _17456_;
  assign _00327_ = w_enq_i & ~(_17862_);
  assign _17863_ = _17856_ | _17458_;
  assign _00328_ = w_enq_i & ~(_17863_);
  assign _17864_ = _17856_ | _17460_;
  assign _00329_ = w_enq_i & ~(_17864_);
  assign _17865_ = _17856_ | _17464_;
  assign _00331_ = w_enq_i & ~(_17865_);
  assign _17866_ = _17856_ | _17466_;
  assign _00332_ = w_enq_i & ~(_17866_);
  assign _17867_ = _17856_ | _17468_;
  assign _00333_ = w_enq_i & ~(_17867_);
  assign _17868_ = _17856_ | _17470_;
  assign _00334_ = w_enq_i & ~(_17868_);
  assign _17869_ = _17856_ | _17473_;
  assign _00335_ = w_enq_i & ~(_17869_);
  assign _17870_ = _17856_ | _17475_;
  assign _00336_ = w_enq_i & ~(_17870_);
  assign _17871_ = _17856_ | _17477_;
  assign _00337_ = w_enq_i & ~(_17871_);
  assign _17872_ = _17856_ | _17479_;
  assign _00338_ = w_enq_i & ~(_17872_);
  assign _17873_ = _17856_ | _17483_;
  assign _00339_ = w_enq_i & ~(_17873_);
  assign _17874_ = _17856_ | _17485_;
  assign _00340_ = w_enq_i & ~(_17874_);
  assign _17875_ = _17856_ | _17487_;
  assign _00342_ = w_enq_i & ~(_17875_);
  assign _17876_ = _17856_ | _17489_;
  assign _00343_ = w_enq_i & ~(_17876_);
  assign _17877_ = _17856_ | _17492_;
  assign _00344_ = w_enq_i & ~(_17877_);
  assign _17878_ = _17856_ | _17494_;
  assign _00345_ = w_enq_i & ~(_17878_);
  assign _17879_ = _17856_ | _17496_;
  assign _00346_ = w_enq_i & ~(_17879_);
  assign _17880_ = _17856_ | _17498_;
  assign _00347_ = w_enq_i & ~(_17880_);
  assign _17881_ = _17856_ | _17502_;
  assign _00348_ = w_enq_i & ~(_17881_);
  assign _17882_ = _17856_ | _17504_;
  assign _00349_ = w_enq_i & ~(_17882_);
  assign _17883_ = _17856_ | _17506_;
  assign _00350_ = w_enq_i & ~(_17883_);
  assign _17884_ = _17856_ | _17508_;
  assign _00351_ = w_enq_i & ~(_17884_);
  assign _17885_ = _17856_ | _17511_;
  assign _00353_ = w_enq_i & ~(_17885_);
  assign _17886_ = _17856_ | _17513_;
  assign _00354_ = w_enq_i & ~(_17886_);
  assign _17887_ = _17856_ | _17515_;
  assign _00355_ = w_enq_i & ~(_17887_);
  assign _17888_ = _17856_ | _17517_;
  assign _00356_ = w_enq_i & ~(_17888_);
  assign _17889_ = _17755_ | _17621_;
  assign _17890_ = _17889_ | _17438_;
  assign _17891_ = _17890_ | _17437_;
  assign _00357_ = w_enq_i & ~(_17891_);
  assign _17892_ = _17890_ | _17444_;
  assign _00358_ = w_enq_i & ~(_17892_);
  assign _17893_ = _17890_ | _17447_;
  assign _00359_ = w_enq_i & ~(_17893_);
  assign _17894_ = _17890_ | _17450_;
  assign _00360_ = w_enq_i & ~(_17894_);
  assign _17895_ = _17890_ | _17454_;
  assign _00361_ = w_enq_i & ~(_17895_);
  assign _17896_ = _17890_ | _17456_;
  assign _00362_ = w_enq_i & ~(_17896_);
  assign _17897_ = _17890_ | _17458_;
  assign _00364_ = w_enq_i & ~(_17897_);
  assign _17898_ = _17890_ | _17460_;
  assign _00365_ = w_enq_i & ~(_17898_);
  assign _17899_ = _17890_ | _17464_;
  assign _00366_ = w_enq_i & ~(_17899_);
  assign _17900_ = _17890_ | _17466_;
  assign _00367_ = w_enq_i & ~(_17900_);
  assign _17901_ = _17890_ | _17468_;
  assign _00368_ = w_enq_i & ~(_17901_);
  assign _17902_ = _17890_ | _17470_;
  assign _00369_ = w_enq_i & ~(_17902_);
  assign _17903_ = _17890_ | _17473_;
  assign _00370_ = w_enq_i & ~(_17903_);
  assign _17904_ = _17890_ | _17475_;
  assign _00371_ = w_enq_i & ~(_17904_);
  assign _17905_ = _17890_ | _17477_;
  assign _00372_ = w_enq_i & ~(_17905_);
  assign _17906_ = _17890_ | _17479_;
  assign _00373_ = w_enq_i & ~(_17906_);
  assign _17907_ = _17890_ | _17483_;
  assign _00376_ = w_enq_i & ~(_17907_);
  assign _17908_ = _17890_ | _17485_;
  assign _00377_ = w_enq_i & ~(_17908_);
  assign _17909_ = _17890_ | _17487_;
  assign _00378_ = w_enq_i & ~(_17909_);
  assign _17910_ = _17890_ | _17489_;
  assign _00379_ = w_enq_i & ~(_17910_);
  assign _17911_ = _17890_ | _17492_;
  assign _00380_ = w_enq_i & ~(_17911_);
  assign _17912_ = _17890_ | _17494_;
  assign _00381_ = w_enq_i & ~(_17912_);
  assign _17913_ = _17890_ | _17496_;
  assign _00382_ = w_enq_i & ~(_17913_);
  assign _17914_ = _17890_ | _17498_;
  assign _00383_ = w_enq_i & ~(_17914_);
  assign _17915_ = _17890_ | _17502_;
  assign _00384_ = w_enq_i & ~(_17915_);
  assign _17916_ = _17890_ | _17504_;
  assign _00385_ = w_enq_i & ~(_17916_);
  assign _17917_ = _17890_ | _17506_;
  assign _00387_ = w_enq_i & ~(_17917_);
  assign _17918_ = _17890_ | _17508_;
  assign _00388_ = w_enq_i & ~(_17918_);
  assign _17919_ = _17890_ | _17511_;
  assign _00389_ = w_enq_i & ~(_17919_);
  assign _17920_ = _17890_ | _17513_;
  assign _00390_ = w_enq_i & ~(_17920_);
  assign _17921_ = _17890_ | _17515_;
  assign _00391_ = w_enq_i & ~(_17921_);
  assign _17922_ = _17890_ | _17517_;
  assign _00392_ = w_enq_i & ~(_17922_);
  assign _17923_ = _17889_ | _17519_;
  assign _17924_ = _17923_ | _17437_;
  assign _00393_ = w_enq_i & ~(_17924_);
  assign _17925_ = _17923_ | _17444_;
  assign _00394_ = w_enq_i & ~(_17925_);
  assign _17926_ = _17923_ | _17447_;
  assign _00395_ = w_enq_i & ~(_17926_);
  assign _17927_ = _17923_ | _17450_;
  assign _00396_ = w_enq_i & ~(_17927_);
  assign _17928_ = _17923_ | _17454_;
  assign _00398_ = w_enq_i & ~(_17928_);
  assign _17929_ = _17923_ | _17456_;
  assign _00399_ = w_enq_i & ~(_17929_);
  assign _17930_ = _17923_ | _17458_;
  assign _00400_ = w_enq_i & ~(_17930_);
  assign _17931_ = _17923_ | _17460_;
  assign _00401_ = w_enq_i & ~(_17931_);
  assign _17932_ = _17923_ | _17464_;
  assign _00402_ = w_enq_i & ~(_17932_);
  assign _17933_ = _17923_ | _17466_;
  assign _00403_ = w_enq_i & ~(_17933_);
  assign _17934_ = _17923_ | _17468_;
  assign _00404_ = w_enq_i & ~(_17934_);
  assign _17935_ = _17923_ | _17470_;
  assign _00405_ = w_enq_i & ~(_17935_);
  assign _17936_ = _17923_ | _17473_;
  assign _00406_ = w_enq_i & ~(_17936_);
  assign _17937_ = _17923_ | _17475_;
  assign _00407_ = w_enq_i & ~(_17937_);
  assign _17938_ = _17923_ | _17477_;
  assign _00409_ = w_enq_i & ~(_17938_);
  assign _17939_ = _17923_ | _17479_;
  assign _00410_ = w_enq_i & ~(_17939_);
  assign _17940_ = _17923_ | _17483_;
  assign _00411_ = w_enq_i & ~(_17940_);
  assign _17941_ = _17923_ | _17485_;
  assign _00412_ = w_enq_i & ~(_17941_);
  assign _17942_ = _17923_ | _17487_;
  assign _00413_ = w_enq_i & ~(_17942_);
  assign _17943_ = _17923_ | _17489_;
  assign _00414_ = w_enq_i & ~(_17943_);
  assign _17944_ = _17923_ | _17492_;
  assign _00415_ = w_enq_i & ~(_17944_);
  assign _17945_ = _17923_ | _17494_;
  assign _00416_ = w_enq_i & ~(_17945_);
  assign _17946_ = _17923_ | _17496_;
  assign _00417_ = w_enq_i & ~(_17946_);
  assign _17947_ = _17923_ | _17498_;
  assign _00418_ = w_enq_i & ~(_17947_);
  assign _17948_ = _17923_ | _17502_;
  assign _00420_ = w_enq_i & ~(_17948_);
  assign _17949_ = _17923_ | _17504_;
  assign _00421_ = w_enq_i & ~(_17949_);
  assign _17950_ = _17923_ | _17506_;
  assign _00422_ = w_enq_i & ~(_17950_);
  assign _17951_ = _17923_ | _17508_;
  assign _00423_ = w_enq_i & ~(_17951_);
  assign _17952_ = _17923_ | _17511_;
  assign _00424_ = w_enq_i & ~(_17952_);
  assign _17953_ = _17923_ | _17513_;
  assign _00425_ = w_enq_i & ~(_17953_);
  assign _17954_ = _17923_ | _17515_;
  assign _00426_ = w_enq_i & ~(_17954_);
  assign _17955_ = _17923_ | _17517_;
  assign _00427_ = w_enq_i & ~(_17955_);
  assign _17956_ = _17889_ | _17553_;
  assign _17957_ = _17956_ | _17437_;
  assign _00428_ = w_enq_i & ~(_17957_);
  assign _17958_ = _17956_ | _17444_;
  assign _00429_ = w_enq_i & ~(_17958_);
  assign _17959_ = _17956_ | _17447_;
  assign _00431_ = w_enq_i & ~(_17959_);
  assign _17960_ = _17956_ | _17450_;
  assign _00432_ = w_enq_i & ~(_17960_);
  assign _17961_ = _17956_ | _17454_;
  assign _00433_ = w_enq_i & ~(_17961_);
  assign _17962_ = _17956_ | _17456_;
  assign _00434_ = w_enq_i & ~(_17962_);
  assign _17963_ = _17956_ | _17458_;
  assign _00435_ = w_enq_i & ~(_17963_);
  assign _17964_ = _17956_ | _17460_;
  assign _00436_ = w_enq_i & ~(_17964_);
  assign _17965_ = _17956_ | _17464_;
  assign _00437_ = w_enq_i & ~(_17965_);
  assign _17966_ = _17956_ | _17466_;
  assign _00438_ = w_enq_i & ~(_17966_);
  assign _17967_ = _17956_ | _17468_;
  assign _00439_ = w_enq_i & ~(_17967_);
  assign _17968_ = _17956_ | _17470_;
  assign _00440_ = w_enq_i & ~(_17968_);
  assign _17969_ = _17956_ | _17473_;
  assign _00442_ = w_enq_i & ~(_17969_);
  assign _17970_ = _17956_ | _17475_;
  assign _00443_ = w_enq_i & ~(_17970_);
  assign _17971_ = _17956_ | _17477_;
  assign _00444_ = w_enq_i & ~(_17971_);
  assign _17972_ = _17956_ | _17479_;
  assign _00445_ = w_enq_i & ~(_17972_);
  assign _17973_ = _17956_ | _17483_;
  assign _00446_ = w_enq_i & ~(_17973_);
  assign _17974_ = _17956_ | _17485_;
  assign _00447_ = w_enq_i & ~(_17974_);
  assign _17975_ = _17956_ | _17487_;
  assign _00448_ = w_enq_i & ~(_17975_);
  assign _17976_ = _17956_ | _17489_;
  assign _00449_ = w_enq_i & ~(_17976_);
  assign _17977_ = _17956_ | _17492_;
  assign _00450_ = w_enq_i & ~(_17977_);
  assign _17978_ = _17956_ | _17494_;
  assign _00451_ = w_enq_i & ~(_17978_);
  assign _17979_ = _17956_ | _17496_;
  assign _00453_ = w_enq_i & ~(_17979_);
  assign _17980_ = _17956_ | _17498_;
  assign _00454_ = w_enq_i & ~(_17980_);
  assign _17981_ = _17956_ | _17502_;
  assign _00455_ = w_enq_i & ~(_17981_);
  assign _17982_ = _17956_ | _17504_;
  assign _00456_ = w_enq_i & ~(_17982_);
  assign _17983_ = _17956_ | _17506_;
  assign _00457_ = w_enq_i & ~(_17983_);
  assign _17984_ = _17956_ | _17508_;
  assign _00458_ = w_enq_i & ~(_17984_);
  assign _17985_ = _17956_ | _17511_;
  assign _00459_ = w_enq_i & ~(_17985_);
  assign _17986_ = _17956_ | _17513_;
  assign _00460_ = w_enq_i & ~(_17986_);
  assign _17987_ = _17956_ | _17515_;
  assign _00461_ = w_enq_i & ~(_17987_);
  assign _17988_ = _17956_ | _17517_;
  assign _00462_ = w_enq_i & ~(_17988_);
  assign _17989_ = _17889_ | _17587_;
  assign _17990_ = _17989_ | _17437_;
  assign _00464_ = w_enq_i & ~(_17990_);
  assign _17991_ = _17989_ | _17444_;
  assign _00465_ = w_enq_i & ~(_17991_);
  assign _17992_ = _17989_ | _17447_;
  assign _00466_ = w_enq_i & ~(_17992_);
  assign _17993_ = _17989_ | _17450_;
  assign _00467_ = w_enq_i & ~(_17993_);
  assign _17994_ = _17989_ | _17454_;
  assign _00468_ = w_enq_i & ~(_17994_);
  assign _17995_ = _17989_ | _17456_;
  assign _00469_ = w_enq_i & ~(_17995_);
  assign _17996_ = _17989_ | _17458_;
  assign _00470_ = w_enq_i & ~(_17996_);
  assign _17997_ = _17989_ | _17460_;
  assign _00471_ = w_enq_i & ~(_17997_);
  assign _17998_ = _17989_ | _17464_;
  assign _00472_ = w_enq_i & ~(_17998_);
  assign _17999_ = _17989_ | _17466_;
  assign _00473_ = w_enq_i & ~(_17999_);
  assign _18000_ = _17989_ | _17468_;
  assign _00475_ = w_enq_i & ~(_18000_);
  assign _18001_ = _17989_ | _17470_;
  assign _00476_ = w_enq_i & ~(_18001_);
  assign _18002_ = _17989_ | _17473_;
  assign _00477_ = w_enq_i & ~(_18002_);
  assign _18003_ = _17989_ | _17475_;
  assign _00478_ = w_enq_i & ~(_18003_);
  assign _18004_ = _17989_ | _17477_;
  assign _00479_ = w_enq_i & ~(_18004_);
  assign _18005_ = _17989_ | _17479_;
  assign _00480_ = w_enq_i & ~(_18005_);
  assign _18006_ = _17989_ | _17483_;
  assign _00481_ = w_enq_i & ~(_18006_);
  assign _18007_ = _17989_ | _17485_;
  assign _00482_ = w_enq_i & ~(_18007_);
  assign _18008_ = _17989_ | _17487_;
  assign _00483_ = w_enq_i & ~(_18008_);
  assign _18009_ = _17989_ | _17489_;
  assign _00484_ = w_enq_i & ~(_18009_);
  assign _18010_ = _17989_ | _17492_;
  assign _00487_ = w_enq_i & ~(_18010_);
  assign _18011_ = _17989_ | _17494_;
  assign _00488_ = w_enq_i & ~(_18011_);
  assign _18012_ = _17989_ | _17496_;
  assign _00489_ = w_enq_i & ~(_18012_);
  assign _18013_ = _17989_ | _17498_;
  assign _00490_ = w_enq_i & ~(_18013_);
  assign _18014_ = _17989_ | _17502_;
  assign _00491_ = w_enq_i & ~(_18014_);
  assign _18015_ = _17989_ | _17504_;
  assign _00492_ = w_enq_i & ~(_18015_);
  assign _18016_ = _17989_ | _17506_;
  assign _00493_ = w_enq_i & ~(_18016_);
  assign _18017_ = _17989_ | _17508_;
  assign _00494_ = w_enq_i & ~(_18017_);
  assign _18018_ = _17989_ | _17511_;
  assign _00495_ = w_enq_i & ~(_18018_);
  assign _18019_ = _17989_ | _17513_;
  assign _00496_ = w_enq_i & ~(_18019_);
  assign _18020_ = _17989_ | _17515_;
  assign _00498_ = w_enq_i & ~(_18020_);
  assign _18021_ = _17989_ | _17517_;
  assign _00499_ = w_enq_i & ~(_18021_);
  assign _18022_ = \bapg_wr.w_ptr_r [8] | ~(\bapg_wr.w_ptr_r [9]);
  assign _18023_ = _18022_ | \bapg_wr.w_ptr_r [7];
  assign _18024_ = _18023_ | _17438_;
  assign _18025_ = _18024_ | _17437_;
  assign _00500_ = w_enq_i & ~(_18025_);
  assign _18026_ = _18024_ | _17444_;
  assign _00501_ = w_enq_i & ~(_18026_);
  assign _18027_ = _18024_ | _17447_;
  assign _00502_ = w_enq_i & ~(_18027_);
  assign _18028_ = _18024_ | _17450_;
  assign _00503_ = w_enq_i & ~(_18028_);
  assign _18029_ = _18024_ | _17454_;
  assign _00504_ = w_enq_i & ~(_18029_);
  assign _18030_ = _18024_ | _17456_;
  assign _00505_ = w_enq_i & ~(_18030_);
  assign _18031_ = _18024_ | _17458_;
  assign _00506_ = w_enq_i & ~(_18031_);
  assign _18032_ = _18024_ | _17460_;
  assign _00507_ = w_enq_i & ~(_18032_);
  assign _18033_ = _18024_ | _17464_;
  assign _00509_ = w_enq_i & ~(_18033_);
  assign _18034_ = _18024_ | _17466_;
  assign _00510_ = w_enq_i & ~(_18034_);
  assign _18035_ = _18024_ | _17468_;
  assign _00511_ = w_enq_i & ~(_18035_);
  assign _18036_ = _18024_ | _17470_;
  assign _00512_ = w_enq_i & ~(_18036_);
  assign _18037_ = _18024_ | _17473_;
  assign _00513_ = w_enq_i & ~(_18037_);
  assign _18038_ = _18024_ | _17475_;
  assign _00514_ = w_enq_i & ~(_18038_);
  assign _18039_ = _18024_ | _17477_;
  assign _00515_ = w_enq_i & ~(_18039_);
  assign _18040_ = _18024_ | _17479_;
  assign _00516_ = w_enq_i & ~(_18040_);
  assign _18041_ = _18024_ | _17483_;
  assign _00517_ = w_enq_i & ~(_18041_);
  assign _18042_ = _18024_ | _17485_;
  assign _00518_ = w_enq_i & ~(_18042_);
  assign _18043_ = _18024_ | _17487_;
  assign _00520_ = w_enq_i & ~(_18043_);
  assign _18044_ = _18024_ | _17489_;
  assign _00521_ = w_enq_i & ~(_18044_);
  assign _18045_ = _18024_ | _17492_;
  assign _00522_ = w_enq_i & ~(_18045_);
  assign _18046_ = _18024_ | _17494_;
  assign _00523_ = w_enq_i & ~(_18046_);
  assign _18047_ = _18024_ | _17496_;
  assign _00524_ = w_enq_i & ~(_18047_);
  assign _18048_ = _18024_ | _17498_;
  assign _00525_ = w_enq_i & ~(_18048_);
  assign _18049_ = _18024_ | _17502_;
  assign _00526_ = w_enq_i & ~(_18049_);
  assign _18050_ = _18024_ | _17504_;
  assign _00527_ = w_enq_i & ~(_18050_);
  assign _18051_ = _18024_ | _17506_;
  assign _00528_ = w_enq_i & ~(_18051_);
  assign _18052_ = _18024_ | _17508_;
  assign _00529_ = w_enq_i & ~(_18052_);
  assign _18053_ = _18024_ | _17511_;
  assign _00531_ = w_enq_i & ~(_18053_);
  assign _18054_ = _18024_ | _17513_;
  assign _00532_ = w_enq_i & ~(_18054_);
  assign _18055_ = _18024_ | _17515_;
  assign _00533_ = w_enq_i & ~(_18055_);
  assign _18056_ = _18024_ | _17517_;
  assign _00534_ = w_enq_i & ~(_18056_);
  assign _18057_ = _18023_ | _17519_;
  assign _18058_ = _18057_ | _17437_;
  assign _00535_ = w_enq_i & ~(_18058_);
  assign _18059_ = _18057_ | _17444_;
  assign _00536_ = w_enq_i & ~(_18059_);
  assign _18060_ = _18057_ | _17447_;
  assign _00537_ = w_enq_i & ~(_18060_);
  assign _18061_ = _18057_ | _17450_;
  assign _00538_ = w_enq_i & ~(_18061_);
  assign _18062_ = _18057_ | _17454_;
  assign _00539_ = w_enq_i & ~(_18062_);
  assign _18063_ = _18057_ | _17456_;
  assign _00540_ = w_enq_i & ~(_18063_);
  assign _18064_ = _18057_ | _17458_;
  assign _00542_ = w_enq_i & ~(_18064_);
  assign _18065_ = _18057_ | _17460_;
  assign _00543_ = w_enq_i & ~(_18065_);
  assign _18066_ = _18057_ | _17464_;
  assign _00544_ = w_enq_i & ~(_18066_);
  assign _18067_ = _18057_ | _17466_;
  assign _00545_ = w_enq_i & ~(_18067_);
  assign _18068_ = _18057_ | _17468_;
  assign _00546_ = w_enq_i & ~(_18068_);
  assign _18069_ = _18057_ | _17470_;
  assign _00547_ = w_enq_i & ~(_18069_);
  assign _18070_ = _18057_ | _17473_;
  assign _00548_ = w_enq_i & ~(_18070_);
  assign _18071_ = _18057_ | _17475_;
  assign _00549_ = w_enq_i & ~(_18071_);
  assign _18072_ = _18057_ | _17477_;
  assign _00550_ = w_enq_i & ~(_18072_);
  assign _18073_ = _18057_ | _17479_;
  assign _00551_ = w_enq_i & ~(_18073_);
  assign _18074_ = _18057_ | _17483_;
  assign _00553_ = w_enq_i & ~(_18074_);
  assign _18075_ = _18057_ | _17485_;
  assign _00554_ = w_enq_i & ~(_18075_);
  assign _18076_ = _18057_ | _17487_;
  assign _00555_ = w_enq_i & ~(_18076_);
  assign _18077_ = _18057_ | _17489_;
  assign _00556_ = w_enq_i & ~(_18077_);
  assign _18078_ = _18057_ | _17492_;
  assign _00557_ = w_enq_i & ~(_18078_);
  assign _18079_ = _18057_ | _17494_;
  assign _00558_ = w_enq_i & ~(_18079_);
  assign _18080_ = _18057_ | _17496_;
  assign _00559_ = w_enq_i & ~(_18080_);
  assign _18081_ = _18057_ | _17498_;
  assign _00560_ = w_enq_i & ~(_18081_);
  assign _18082_ = _18057_ | _17502_;
  assign _00561_ = w_enq_i & ~(_18082_);
  assign _18083_ = _18057_ | _17504_;
  assign _00562_ = w_enq_i & ~(_18083_);
  assign _18084_ = _18057_ | _17506_;
  assign _00564_ = w_enq_i & ~(_18084_);
  assign _18085_ = _18057_ | _17508_;
  assign _00565_ = w_enq_i & ~(_18085_);
  assign _18086_ = _18057_ | _17511_;
  assign _00566_ = w_enq_i & ~(_18086_);
  assign _18087_ = _18057_ | _17513_;
  assign _00567_ = w_enq_i & ~(_18087_);
  assign _18088_ = _18057_ | _17515_;
  assign _00568_ = w_enq_i & ~(_18088_);
  assign _18089_ = _18057_ | _17517_;
  assign _00569_ = w_enq_i & ~(_18089_);
  assign _18090_ = _18023_ | _17553_;
  assign _18091_ = _18090_ | _17437_;
  assign _00570_ = w_enq_i & ~(_18091_);
  assign _18092_ = _18090_ | _17444_;
  assign _00571_ = w_enq_i & ~(_18092_);
  assign _18093_ = _18090_ | _17447_;
  assign _00572_ = w_enq_i & ~(_18093_);
  assign _18094_ = _18090_ | _17450_;
  assign _00573_ = w_enq_i & ~(_18094_);
  assign _18095_ = _18090_ | _17454_;
  assign _00575_ = w_enq_i & ~(_18095_);
  assign _18096_ = _18090_ | _17456_;
  assign _00576_ = w_enq_i & ~(_18096_);
  assign _18097_ = _18090_ | _17458_;
  assign _00577_ = w_enq_i & ~(_18097_);
  assign _18098_ = _18090_ | _17460_;
  assign _00578_ = w_enq_i & ~(_18098_);
  assign _18099_ = _18090_ | _17464_;
  assign _00579_ = w_enq_i & ~(_18099_);
  assign _18100_ = _18090_ | _17466_;
  assign _00580_ = w_enq_i & ~(_18100_);
  assign _18101_ = _18090_ | _17468_;
  assign _00581_ = w_enq_i & ~(_18101_);
  assign _18102_ = _18090_ | _17470_;
  assign _00582_ = w_enq_i & ~(_18102_);
  assign _18103_ = _18090_ | _17473_;
  assign _00583_ = w_enq_i & ~(_18103_);
  assign _18104_ = _18090_ | _17475_;
  assign _00584_ = w_enq_i & ~(_18104_);
  assign _18105_ = _18090_ | _17477_;
  assign _00586_ = w_enq_i & ~(_18105_);
  assign _18106_ = _18090_ | _17479_;
  assign _00587_ = w_enq_i & ~(_18106_);
  assign _18107_ = _18090_ | _17483_;
  assign _00588_ = w_enq_i & ~(_18107_);
  assign _18108_ = _18090_ | _17485_;
  assign _00589_ = w_enq_i & ~(_18108_);
  assign _18109_ = _18090_ | _17487_;
  assign _00590_ = w_enq_i & ~(_18109_);
  assign _18110_ = _18090_ | _17489_;
  assign _00591_ = w_enq_i & ~(_18110_);
  assign _18111_ = _18090_ | _17492_;
  assign _00592_ = w_enq_i & ~(_18111_);
  assign _18112_ = _18090_ | _17494_;
  assign _00593_ = w_enq_i & ~(_18112_);
  assign _18113_ = _18090_ | _17496_;
  assign _00594_ = w_enq_i & ~(_18113_);
  assign _18114_ = _18090_ | _17498_;
  assign _00595_ = w_enq_i & ~(_18114_);
  assign _18115_ = _18090_ | _17502_;
  assign _00598_ = w_enq_i & ~(_18115_);
  assign _18116_ = _18090_ | _17504_;
  assign _00599_ = w_enq_i & ~(_18116_);
  assign _18117_ = _18090_ | _17506_;
  assign _00600_ = w_enq_i & ~(_18117_);
  assign _18118_ = _18090_ | _17508_;
  assign _00601_ = w_enq_i & ~(_18118_);
  assign _18119_ = _18090_ | _17511_;
  assign _00602_ = w_enq_i & ~(_18119_);
  assign _18120_ = _18090_ | _17513_;
  assign _00603_ = w_enq_i & ~(_18120_);
  assign _18121_ = _18090_ | _17515_;
  assign _00604_ = w_enq_i & ~(_18121_);
  assign _18122_ = _18090_ | _17517_;
  assign _00605_ = w_enq_i & ~(_18122_);
  assign _18123_ = _18023_ | _17587_;
  assign _18124_ = _18123_ | _17437_;
  assign _00606_ = w_enq_i & ~(_18124_);
  assign _18125_ = _18123_ | _17444_;
  assign _00607_ = w_enq_i & ~(_18125_);
  assign _18126_ = _18123_ | _17447_;
  assign _00609_ = w_enq_i & ~(_18126_);
  assign _18127_ = _18123_ | _17450_;
  assign _00610_ = w_enq_i & ~(_18127_);
  assign _18128_ = _18123_ | _17454_;
  assign _00611_ = w_enq_i & ~(_18128_);
  assign _18129_ = _18123_ | _17456_;
  assign _00612_ = w_enq_i & ~(_18129_);
  assign _18130_ = _18123_ | _17458_;
  assign _00613_ = w_enq_i & ~(_18130_);
  assign _18131_ = _18123_ | _17460_;
  assign _00614_ = w_enq_i & ~(_18131_);
  assign _18132_ = _18123_ | _17464_;
  assign _00615_ = w_enq_i & ~(_18132_);
  assign _18133_ = _18123_ | _17466_;
  assign _00616_ = w_enq_i & ~(_18133_);
  assign _18134_ = _18123_ | _17468_;
  assign _00617_ = w_enq_i & ~(_18134_);
  assign _18135_ = _18123_ | _17470_;
  assign _00618_ = w_enq_i & ~(_18135_);
  assign _18136_ = _18123_ | _17473_;
  assign _00620_ = w_enq_i & ~(_18136_);
  assign _18137_ = _18123_ | _17475_;
  assign _00621_ = w_enq_i & ~(_18137_);
  assign _18138_ = _18123_ | _17477_;
  assign _00622_ = w_enq_i & ~(_18138_);
  assign _18139_ = _18123_ | _17479_;
  assign _00623_ = w_enq_i & ~(_18139_);
  assign _18140_ = _18123_ | _17483_;
  assign _00624_ = w_enq_i & ~(_18140_);
  assign _18141_ = _18123_ | _17485_;
  assign _00625_ = w_enq_i & ~(_18141_);
  assign _18142_ = _18123_ | _17487_;
  assign _00626_ = w_enq_i & ~(_18142_);
  assign _18143_ = _18123_ | _17489_;
  assign _00627_ = w_enq_i & ~(_18143_);
  assign _18144_ = _18123_ | _17492_;
  assign _00628_ = w_enq_i & ~(_18144_);
  assign _18145_ = _18123_ | _17494_;
  assign _00629_ = w_enq_i & ~(_18145_);
  assign _18146_ = _18123_ | _17496_;
  assign _00631_ = w_enq_i & ~(_18146_);
  assign _18147_ = _18123_ | _17498_;
  assign _00632_ = w_enq_i & ~(_18147_);
  assign _18148_ = _18123_ | _17502_;
  assign _00633_ = w_enq_i & ~(_18148_);
  assign _18149_ = _18123_ | _17504_;
  assign _00634_ = w_enq_i & ~(_18149_);
  assign _18150_ = _18123_ | _17506_;
  assign _00635_ = w_enq_i & ~(_18150_);
  assign _18151_ = _18123_ | _17508_;
  assign _00636_ = w_enq_i & ~(_18151_);
  assign _18152_ = _18123_ | _17511_;
  assign _00637_ = w_enq_i & ~(_18152_);
  assign _18153_ = _18123_ | _17513_;
  assign _00638_ = w_enq_i & ~(_18153_);
  assign _18154_ = _18123_ | _17515_;
  assign _00639_ = w_enq_i & ~(_18154_);
  assign _18155_ = _18123_ | _17517_;
  assign _00640_ = w_enq_i & ~(_18155_);
  assign _18156_ = _18022_ | _17621_;
  assign _18157_ = _18156_ | _17438_;
  assign _18158_ = _18157_ | _17437_;
  assign _00642_ = w_enq_i & ~(_18158_);
  assign _18159_ = _18157_ | _17444_;
  assign _00643_ = w_enq_i & ~(_18159_);
  assign _18160_ = _18157_ | _17447_;
  assign _00644_ = w_enq_i & ~(_18160_);
  assign _18161_ = _18157_ | _17450_;
  assign _00645_ = w_enq_i & ~(_18161_);
  assign _18162_ = _18157_ | _17454_;
  assign _00646_ = w_enq_i & ~(_18162_);
  assign _18163_ = _18157_ | _17456_;
  assign _00647_ = w_enq_i & ~(_18163_);
  assign _18164_ = _18157_ | _17458_;
  assign _00648_ = w_enq_i & ~(_18164_);
  assign _18165_ = _18157_ | _17460_;
  assign _00649_ = w_enq_i & ~(_18165_);
  assign _18166_ = _18157_ | _17464_;
  assign _00650_ = w_enq_i & ~(_18166_);
  assign _18167_ = _18157_ | _17466_;
  assign _00651_ = w_enq_i & ~(_18167_);
  assign _18168_ = _18157_ | _17468_;
  assign _00653_ = w_enq_i & ~(_18168_);
  assign _18169_ = _18157_ | _17470_;
  assign _00654_ = w_enq_i & ~(_18169_);
  assign _18170_ = _18157_ | _17473_;
  assign _00655_ = w_enq_i & ~(_18170_);
  assign _18171_ = _18157_ | _17475_;
  assign _00656_ = w_enq_i & ~(_18171_);
  assign _18172_ = _18157_ | _17477_;
  assign _00657_ = w_enq_i & ~(_18172_);
  assign _18173_ = _18157_ | _17479_;
  assign _00658_ = w_enq_i & ~(_18173_);
  assign _18174_ = _18157_ | _17483_;
  assign _00659_ = w_enq_i & ~(_18174_);
  assign _18175_ = _18157_ | _17485_;
  assign _00660_ = w_enq_i & ~(_18175_);
  assign _18176_ = _18157_ | _17487_;
  assign _00661_ = w_enq_i & ~(_18176_);
  assign _18177_ = _18157_ | _17489_;
  assign _00662_ = w_enq_i & ~(_18177_);
  assign _18178_ = _18157_ | _17492_;
  assign _00664_ = w_enq_i & ~(_18178_);
  assign _18179_ = _18157_ | _17494_;
  assign _00665_ = w_enq_i & ~(_18179_);
  assign _18180_ = _18157_ | _17496_;
  assign _00666_ = w_enq_i & ~(_18180_);
  assign _18181_ = _18157_ | _17498_;
  assign _00667_ = w_enq_i & ~(_18181_);
  assign _18182_ = _18157_ | _17502_;
  assign _00668_ = w_enq_i & ~(_18182_);
  assign _18183_ = _18157_ | _17504_;
  assign _00669_ = w_enq_i & ~(_18183_);
  assign _18184_ = _18157_ | _17506_;
  assign _00670_ = w_enq_i & ~(_18184_);
  assign _18185_ = _18157_ | _17508_;
  assign _00671_ = w_enq_i & ~(_18185_);
  assign _18186_ = _18157_ | _17511_;
  assign _00672_ = w_enq_i & ~(_18186_);
  assign _18187_ = _18157_ | _17513_;
  assign _00673_ = w_enq_i & ~(_18187_);
  assign _18188_ = _18157_ | _17515_;
  assign _00675_ = w_enq_i & ~(_18188_);
  assign _18189_ = _18157_ | _17517_;
  assign _00676_ = w_enq_i & ~(_18189_);
  assign _18190_ = _18156_ | _17519_;
  assign _18191_ = _18190_ | _17437_;
  assign _00677_ = w_enq_i & ~(_18191_);
  assign _18192_ = _18190_ | _17444_;
  assign _00678_ = w_enq_i & ~(_18192_);
  assign _18193_ = _18190_ | _17447_;
  assign _00679_ = w_enq_i & ~(_18193_);
  assign _18194_ = _18190_ | _17450_;
  assign _00680_ = w_enq_i & ~(_18194_);
  assign _18195_ = _18190_ | _17454_;
  assign _00681_ = w_enq_i & ~(_18195_);
  assign _18196_ = _18190_ | _17456_;
  assign _00682_ = w_enq_i & ~(_18196_);
  assign _18197_ = _18190_ | _17458_;
  assign _00683_ = w_enq_i & ~(_18197_);
  assign _18198_ = _18190_ | _17460_;
  assign _00684_ = w_enq_i & ~(_18198_);
  assign _18199_ = _18190_ | _17464_;
  assign _00686_ = w_enq_i & ~(_18199_);
  assign _18200_ = _18190_ | _17466_;
  assign _00687_ = w_enq_i & ~(_18200_);
  assign _18201_ = _18190_ | _17468_;
  assign _00688_ = w_enq_i & ~(_18201_);
  assign _18202_ = _18190_ | _17470_;
  assign _00689_ = w_enq_i & ~(_18202_);
  assign _18203_ = _18190_ | _17473_;
  assign _00690_ = w_enq_i & ~(_18203_);
  assign _18204_ = _18190_ | _17475_;
  assign _00691_ = w_enq_i & ~(_18204_);
  assign _18205_ = _18190_ | _17477_;
  assign _00692_ = w_enq_i & ~(_18205_);
  assign _18206_ = _18190_ | _17479_;
  assign _00693_ = w_enq_i & ~(_18206_);
  assign _18207_ = _18190_ | _17483_;
  assign _00694_ = w_enq_i & ~(_18207_);
  assign _18208_ = _18190_ | _17485_;
  assign _00695_ = w_enq_i & ~(_18208_);
  assign _18209_ = _18190_ | _17487_;
  assign _00697_ = w_enq_i & ~(_18209_);
  assign _18210_ = _18190_ | _17489_;
  assign _00698_ = w_enq_i & ~(_18210_);
  assign _18211_ = _18190_ | _17492_;
  assign _00699_ = w_enq_i & ~(_18211_);
  assign _18212_ = _18190_ | _17494_;
  assign _00700_ = w_enq_i & ~(_18212_);
  assign _18213_ = _18190_ | _17496_;
  assign _00701_ = w_enq_i & ~(_18213_);
  assign _18214_ = _18190_ | _17498_;
  assign _00702_ = w_enq_i & ~(_18214_);
  assign _18215_ = _18190_ | _17502_;
  assign _00703_ = w_enq_i & ~(_18215_);
  assign _18216_ = _18190_ | _17504_;
  assign _00704_ = w_enq_i & ~(_18216_);
  assign _18217_ = _18190_ | _17506_;
  assign _00705_ = w_enq_i & ~(_18217_);
  assign _18218_ = _18190_ | _17508_;
  assign _00706_ = w_enq_i & ~(_18218_);
  assign _18219_ = _18190_ | _17511_;
  assign _00709_ = w_enq_i & ~(_18219_);
  assign _18220_ = _18190_ | _17513_;
  assign _00710_ = w_enq_i & ~(_18220_);
  assign _18221_ = _18190_ | _17515_;
  assign _00711_ = w_enq_i & ~(_18221_);
  assign _18222_ = _18190_ | _17517_;
  assign _00712_ = w_enq_i & ~(_18222_);
  assign _18223_ = _18156_ | _17553_;
  assign _18224_ = _18223_ | _17437_;
  assign _00713_ = w_enq_i & ~(_18224_);
  assign _18225_ = _18223_ | _17444_;
  assign _00714_ = w_enq_i & ~(_18225_);
  assign _18226_ = _18223_ | _17447_;
  assign _00715_ = w_enq_i & ~(_18226_);
  assign _18227_ = _18223_ | _17450_;
  assign _00716_ = w_enq_i & ~(_18227_);
  assign _18228_ = _18223_ | _17454_;
  assign _00717_ = w_enq_i & ~(_18228_);
  assign _18229_ = _18223_ | _17456_;
  assign _00718_ = w_enq_i & ~(_18229_);
  assign _18230_ = _18223_ | _17458_;
  assign _00720_ = w_enq_i & ~(_18230_);
  assign _18231_ = _18223_ | _17460_;
  assign _00721_ = w_enq_i & ~(_18231_);
  assign _18232_ = _18223_ | _17464_;
  assign _00722_ = w_enq_i & ~(_18232_);
  assign _18233_ = _18223_ | _17466_;
  assign _00723_ = w_enq_i & ~(_18233_);
  assign _18234_ = _18223_ | _17468_;
  assign _00724_ = w_enq_i & ~(_18234_);
  assign _18235_ = _18223_ | _17470_;
  assign _00725_ = w_enq_i & ~(_18235_);
  assign _18236_ = _18223_ | _17473_;
  assign _00726_ = w_enq_i & ~(_18236_);
  assign _18237_ = _18223_ | _17475_;
  assign _00727_ = w_enq_i & ~(_18237_);
  assign _18238_ = _18223_ | _17477_;
  assign _00728_ = w_enq_i & ~(_18238_);
  assign _18239_ = _18223_ | _17479_;
  assign _00729_ = w_enq_i & ~(_18239_);
  assign _18240_ = _18223_ | _17483_;
  assign _00731_ = w_enq_i & ~(_18240_);
  assign _18241_ = _18223_ | _17485_;
  assign _00732_ = w_enq_i & ~(_18241_);
  assign _18242_ = _18223_ | _17487_;
  assign _00733_ = w_enq_i & ~(_18242_);
  assign _18243_ = _18223_ | _17489_;
  assign _00734_ = w_enq_i & ~(_18243_);
  assign _18244_ = _18223_ | _17492_;
  assign _00735_ = w_enq_i & ~(_18244_);
  assign _18245_ = _18223_ | _17494_;
  assign _00736_ = w_enq_i & ~(_18245_);
  assign _18246_ = _18223_ | _17496_;
  assign _00737_ = w_enq_i & ~(_18246_);
  assign _18247_ = _18223_ | _17498_;
  assign _00738_ = w_enq_i & ~(_18247_);
  assign _18248_ = _18223_ | _17502_;
  assign _00739_ = w_enq_i & ~(_18248_);
  assign _18249_ = _18223_ | _17504_;
  assign _00740_ = w_enq_i & ~(_18249_);
  assign _18250_ = _18223_ | _17506_;
  assign _00742_ = w_enq_i & ~(_18250_);
  assign _18251_ = _18223_ | _17508_;
  assign _00743_ = w_enq_i & ~(_18251_);
  assign _18252_ = _18223_ | _17511_;
  assign _00744_ = w_enq_i & ~(_18252_);
  assign _18253_ = _18223_ | _17513_;
  assign _00745_ = w_enq_i & ~(_18253_);
  assign _18254_ = _18223_ | _17515_;
  assign _00746_ = w_enq_i & ~(_18254_);
  assign _18255_ = _18223_ | _17517_;
  assign _00747_ = w_enq_i & ~(_18255_);
  assign _18256_ = _18156_ | _17587_;
  assign _18257_ = _18256_ | _17437_;
  assign _00748_ = w_enq_i & ~(_18257_);
  assign _18258_ = _18256_ | _17444_;
  assign _00749_ = w_enq_i & ~(_18258_);
  assign _18259_ = _18256_ | _17447_;
  assign _00750_ = w_enq_i & ~(_18259_);
  assign _18260_ = _18256_ | _17450_;
  assign _00751_ = w_enq_i & ~(_18260_);
  assign _18261_ = _18256_ | _17454_;
  assign _00753_ = w_enq_i & ~(_18261_);
  assign _18262_ = _18256_ | _17456_;
  assign _00754_ = w_enq_i & ~(_18262_);
  assign _18263_ = _18256_ | _17458_;
  assign _00755_ = w_enq_i & ~(_18263_);
  assign _18264_ = _18256_ | _17460_;
  assign _00756_ = w_enq_i & ~(_18264_);
  assign _18265_ = _18256_ | _17464_;
  assign _00757_ = w_enq_i & ~(_18265_);
  assign _18266_ = _18256_ | _17466_;
  assign _00758_ = w_enq_i & ~(_18266_);
  assign _18267_ = _18256_ | _17468_;
  assign _00759_ = w_enq_i & ~(_18267_);
  assign _18268_ = _18256_ | _17470_;
  assign _00760_ = w_enq_i & ~(_18268_);
  assign _18269_ = _18256_ | _17473_;
  assign _00761_ = w_enq_i & ~(_18269_);
  assign _18270_ = _18256_ | _17475_;
  assign _00762_ = w_enq_i & ~(_18270_);
  assign _18271_ = _18256_ | _17477_;
  assign _00764_ = w_enq_i & ~(_18271_);
  assign _18272_ = _18256_ | _17479_;
  assign _00765_ = w_enq_i & ~(_18272_);
  assign _18273_ = _18256_ | _17483_;
  assign _00766_ = w_enq_i & ~(_18273_);
  assign _18274_ = _18256_ | _17485_;
  assign _00767_ = w_enq_i & ~(_18274_);
  assign _18275_ = _18256_ | _17487_;
  assign _00768_ = w_enq_i & ~(_18275_);
  assign _18276_ = _18256_ | _17489_;
  assign _00769_ = w_enq_i & ~(_18276_);
  assign _18277_ = _18256_ | _17492_;
  assign _00770_ = w_enq_i & ~(_18277_);
  assign _18278_ = _18256_ | _17494_;
  assign _00771_ = w_enq_i & ~(_18278_);
  assign _18279_ = _18256_ | _17496_;
  assign _00772_ = w_enq_i & ~(_18279_);
  assign _18280_ = _18256_ | _17498_;
  assign _00773_ = w_enq_i & ~(_18280_);
  assign _18281_ = _18256_ | _17502_;
  assign _00775_ = w_enq_i & ~(_18281_);
  assign _18282_ = _18256_ | _17504_;
  assign _00776_ = w_enq_i & ~(_18282_);
  assign _18283_ = _18256_ | _17506_;
  assign _00777_ = w_enq_i & ~(_18283_);
  assign _18284_ = _18256_ | _17508_;
  assign _00778_ = w_enq_i & ~(_18284_);
  assign _18285_ = _18256_ | _17511_;
  assign _00779_ = w_enq_i & ~(_18285_);
  assign _18286_ = _18256_ | _17513_;
  assign _00780_ = w_enq_i & ~(_18286_);
  assign _18287_ = _18256_ | _17515_;
  assign _00781_ = w_enq_i & ~(_18287_);
  assign _18288_ = _18256_ | _17517_;
  assign _00782_ = w_enq_i & ~(_18288_);
  assign _18289_ = ~(\bapg_wr.w_ptr_r [9] & \bapg_wr.w_ptr_r [8]);
  assign _18290_ = _18289_ | \bapg_wr.w_ptr_r [7];
  assign _18291_ = _18290_ | _17438_;
  assign _18292_ = _18291_ | _17437_;
  assign _00783_ = w_enq_i & ~(_18292_);
  assign _18293_ = _18291_ | _17444_;
  assign _00784_ = w_enq_i & ~(_18293_);
  assign _18294_ = _18291_ | _17447_;
  assign _00786_ = w_enq_i & ~(_18294_);
  assign _18295_ = _18291_ | _17450_;
  assign _00787_ = w_enq_i & ~(_18295_);
  assign _18296_ = _18291_ | _17454_;
  assign _00788_ = w_enq_i & ~(_18296_);
  assign _18297_ = _18291_ | _17456_;
  assign _00789_ = w_enq_i & ~(_18297_);
  assign _18298_ = _18291_ | _17458_;
  assign _00790_ = w_enq_i & ~(_18298_);
  assign _18299_ = _18291_ | _17460_;
  assign _00791_ = w_enq_i & ~(_18299_);
  assign _18300_ = _18291_ | _17464_;
  assign _00792_ = w_enq_i & ~(_18300_);
  assign _18301_ = _18291_ | _17466_;
  assign _00793_ = w_enq_i & ~(_18301_);
  assign _18302_ = _18291_ | _17468_;
  assign _00794_ = w_enq_i & ~(_18302_);
  assign _18303_ = _18291_ | _17470_;
  assign _00795_ = w_enq_i & ~(_18303_);
  assign _18304_ = _18291_ | _17473_;
  assign _00797_ = w_enq_i & ~(_18304_);
  assign _18305_ = _18291_ | _17475_;
  assign _00798_ = w_enq_i & ~(_18305_);
  assign _18306_ = _18291_ | _17477_;
  assign _00799_ = w_enq_i & ~(_18306_);
  assign _18307_ = _18291_ | _17479_;
  assign _00800_ = w_enq_i & ~(_18307_);
  assign _18308_ = _18291_ | _17483_;
  assign _00801_ = w_enq_i & ~(_18308_);
  assign _18309_ = _18291_ | _17485_;
  assign _00802_ = w_enq_i & ~(_18309_);
  assign _18310_ = _18291_ | _17487_;
  assign _00803_ = w_enq_i & ~(_18310_);
  assign _18311_ = _18291_ | _17489_;
  assign _00804_ = w_enq_i & ~(_18311_);
  assign _18312_ = _18291_ | _17492_;
  assign _00805_ = w_enq_i & ~(_18312_);
  assign _18313_ = _18291_ | _17494_;
  assign _00806_ = w_enq_i & ~(_18313_);
  assign _18314_ = _18291_ | _17496_;
  assign _00808_ = w_enq_i & ~(_18314_);
  assign _18315_ = _18291_ | _17498_;
  assign _00809_ = w_enq_i & ~(_18315_);
  assign _18316_ = _18291_ | _17502_;
  assign _00810_ = w_enq_i & ~(_18316_);
  assign _18317_ = _18291_ | _17504_;
  assign _00811_ = w_enq_i & ~(_18317_);
  assign _18318_ = _18291_ | _17506_;
  assign _00812_ = w_enq_i & ~(_18318_);
  assign _18319_ = _18291_ | _17508_;
  assign _00813_ = w_enq_i & ~(_18319_);
  assign _18320_ = _18291_ | _17511_;
  assign _00814_ = w_enq_i & ~(_18320_);
  assign _18321_ = _18291_ | _17513_;
  assign _00815_ = w_enq_i & ~(_18321_);
  assign _18322_ = _18291_ | _17515_;
  assign _00816_ = w_enq_i & ~(_18322_);
  assign _18323_ = _18291_ | _17517_;
  assign _00817_ = w_enq_i & ~(_18323_);
  assign _18324_ = _18290_ | _17519_;
  assign _18325_ = _18324_ | _17437_;
  assign _00820_ = w_enq_i & ~(_18325_);
  assign _18326_ = _18324_ | _17444_;
  assign _00821_ = w_enq_i & ~(_18326_);
  assign _18327_ = _18324_ | _17447_;
  assign _00822_ = w_enq_i & ~(_18327_);
  assign _18328_ = _18324_ | _17450_;
  assign _00823_ = w_enq_i & ~(_18328_);
  assign _18329_ = _18324_ | _17454_;
  assign _00824_ = w_enq_i & ~(_18329_);
  assign _18330_ = _18324_ | _17456_;
  assign _00825_ = w_enq_i & ~(_18330_);
  assign _18331_ = _18324_ | _17458_;
  assign _00826_ = w_enq_i & ~(_18331_);
  assign _18332_ = _18324_ | _17460_;
  assign _00827_ = w_enq_i & ~(_18332_);
  assign _18333_ = _18324_ | _17464_;
  assign _00828_ = w_enq_i & ~(_18333_);
  assign _18334_ = _18324_ | _17466_;
  assign _00829_ = w_enq_i & ~(_18334_);
  assign _18335_ = _18324_ | _17468_;
  assign _00831_ = w_enq_i & ~(_18335_);
  assign _18336_ = _18324_ | _17470_;
  assign _00832_ = w_enq_i & ~(_18336_);
  assign _18337_ = _18324_ | _17473_;
  assign _00833_ = w_enq_i & ~(_18337_);
  assign _18338_ = _18324_ | _17475_;
  assign _00834_ = w_enq_i & ~(_18338_);
  assign _18339_ = _18324_ | _17477_;
  assign _00835_ = w_enq_i & ~(_18339_);
  assign _18340_ = _18324_ | _17479_;
  assign _00836_ = w_enq_i & ~(_18340_);
  assign _18341_ = _18324_ | _17483_;
  assign _00837_ = w_enq_i & ~(_18341_);
  assign _18342_ = _18324_ | _17485_;
  assign _00838_ = w_enq_i & ~(_18342_);
  assign _18343_ = _18324_ | _17487_;
  assign _00839_ = w_enq_i & ~(_18343_);
  assign _18344_ = _18324_ | _17489_;
  assign _00840_ = w_enq_i & ~(_18344_);
  assign _18345_ = _18324_ | _17492_;
  assign _00842_ = w_enq_i & ~(_18345_);
  assign _18346_ = _18324_ | _17494_;
  assign _00843_ = w_enq_i & ~(_18346_);
  assign _18347_ = _18324_ | _17496_;
  assign _00844_ = w_enq_i & ~(_18347_);
  assign _18348_ = _18324_ | _17498_;
  assign _00845_ = w_enq_i & ~(_18348_);
  assign _18349_ = _18324_ | _17502_;
  assign _00846_ = w_enq_i & ~(_18349_);
  assign _18350_ = _18324_ | _17504_;
  assign _00847_ = w_enq_i & ~(_18350_);
  assign _18351_ = _18324_ | _17506_;
  assign _00848_ = w_enq_i & ~(_18351_);
  assign _18352_ = _18324_ | _17508_;
  assign _00849_ = w_enq_i & ~(_18352_);
  assign _18353_ = _18324_ | _17511_;
  assign _00850_ = w_enq_i & ~(_18353_);
  assign _18354_ = _18324_ | _17513_;
  assign _00851_ = w_enq_i & ~(_18354_);
  assign _18355_ = _18324_ | _17515_;
  assign _00853_ = w_enq_i & ~(_18355_);
  assign _18356_ = _18324_ | _17517_;
  assign _00854_ = w_enq_i & ~(_18356_);
  assign _18357_ = _18290_ | _17553_;
  assign _18358_ = _18357_ | _17437_;
  assign _00855_ = w_enq_i & ~(_18358_);
  assign _18359_ = _18357_ | _17444_;
  assign _00856_ = w_enq_i & ~(_18359_);
  assign _18360_ = _18357_ | _17447_;
  assign _00857_ = w_enq_i & ~(_18360_);
  assign _18361_ = _18357_ | _17450_;
  assign _00858_ = w_enq_i & ~(_18361_);
  assign _18362_ = _18357_ | _17454_;
  assign _00859_ = w_enq_i & ~(_18362_);
  assign _18363_ = _18357_ | _17456_;
  assign _00860_ = w_enq_i & ~(_18363_);
  assign _18364_ = _18357_ | _17458_;
  assign _00861_ = w_enq_i & ~(_18364_);
  assign _18365_ = _18357_ | _17460_;
  assign _00862_ = w_enq_i & ~(_18365_);
  assign _18366_ = _18357_ | _17464_;
  assign _00864_ = w_enq_i & ~(_18366_);
  assign _18367_ = _18357_ | _17466_;
  assign _00865_ = w_enq_i & ~(_18367_);
  assign _18368_ = _18357_ | _17468_;
  assign _00866_ = w_enq_i & ~(_18368_);
  assign _18369_ = _18357_ | _17470_;
  assign _00867_ = w_enq_i & ~(_18369_);
  assign _18370_ = _18357_ | _17473_;
  assign _00868_ = w_enq_i & ~(_18370_);
  assign _18371_ = _18357_ | _17475_;
  assign _00869_ = w_enq_i & ~(_18371_);
  assign _18372_ = _18357_ | _17477_;
  assign _00870_ = w_enq_i & ~(_18372_);
  assign _18373_ = _18357_ | _17479_;
  assign _00871_ = w_enq_i & ~(_18373_);
  assign _18374_ = _18357_ | _17483_;
  assign _00872_ = w_enq_i & ~(_18374_);
  assign _18375_ = _18357_ | _17485_;
  assign _00873_ = w_enq_i & ~(_18375_);
  assign _18376_ = _18357_ | _17487_;
  assign _00875_ = w_enq_i & ~(_18376_);
  assign _18377_ = _18357_ | _17489_;
  assign _00876_ = w_enq_i & ~(_18377_);
  assign _18378_ = _18357_ | _17492_;
  assign _00877_ = w_enq_i & ~(_18378_);
  assign _18379_ = _18357_ | _17494_;
  assign _00878_ = w_enq_i & ~(_18379_);
  assign _18380_ = _18357_ | _17496_;
  assign _00879_ = w_enq_i & ~(_18380_);
  assign _18381_ = _18357_ | _17498_;
  assign _00880_ = w_enq_i & ~(_18381_);
  assign _18382_ = _18357_ | _17502_;
  assign _00881_ = w_enq_i & ~(_18382_);
  assign _18383_ = _18357_ | _17504_;
  assign _00882_ = w_enq_i & ~(_18383_);
  assign _18384_ = _18357_ | _17506_;
  assign _00883_ = w_enq_i & ~(_18384_);
  assign _18385_ = _18357_ | _17508_;
  assign _00884_ = w_enq_i & ~(_18385_);
  assign _18386_ = _18357_ | _17511_;
  assign _00886_ = w_enq_i & ~(_18386_);
  assign _18387_ = _18357_ | _17513_;
  assign _00887_ = w_enq_i & ~(_18387_);
  assign _18388_ = _18357_ | _17515_;
  assign _00888_ = w_enq_i & ~(_18388_);
  assign _18389_ = _18357_ | _17517_;
  assign _00889_ = w_enq_i & ~(_18389_);
  assign _18390_ = _18290_ | _17587_;
  assign _18391_ = _18390_ | _17437_;
  assign _00890_ = w_enq_i & ~(_18391_);
  assign _18392_ = _18390_ | _17444_;
  assign _00891_ = w_enq_i & ~(_18392_);
  assign _18393_ = _18390_ | _17447_;
  assign _00892_ = w_enq_i & ~(_18393_);
  assign _18394_ = _18390_ | _17450_;
  assign _00893_ = w_enq_i & ~(_18394_);
  assign _18395_ = _18390_ | _17454_;
  assign _00894_ = w_enq_i & ~(_18395_);
  assign _18396_ = _18390_ | _17456_;
  assign _00895_ = w_enq_i & ~(_18396_);
  assign _18397_ = _18390_ | _17458_;
  assign _00897_ = w_enq_i & ~(_18397_);
  assign _18398_ = _18390_ | _17460_;
  assign _00898_ = w_enq_i & ~(_18398_);
  assign _18399_ = _18390_ | _17464_;
  assign _00899_ = w_enq_i & ~(_18399_);
  assign _18400_ = _18390_ | _17466_;
  assign _00900_ = w_enq_i & ~(_18400_);
  assign _18401_ = _18390_ | _17468_;
  assign _00901_ = w_enq_i & ~(_18401_);
  assign _18402_ = _18390_ | _17470_;
  assign _00902_ = w_enq_i & ~(_18402_);
  assign _18403_ = _18390_ | _17473_;
  assign _00903_ = w_enq_i & ~(_18403_);
  assign _18404_ = _18390_ | _17475_;
  assign _00904_ = w_enq_i & ~(_18404_);
  assign _18405_ = _18390_ | _17477_;
  assign _00905_ = w_enq_i & ~(_18405_);
  assign _18406_ = _18390_ | _17479_;
  assign _00906_ = w_enq_i & ~(_18406_);
  assign _18407_ = _18390_ | _17483_;
  assign _00908_ = w_enq_i & ~(_18407_);
  assign _18408_ = _18390_ | _17485_;
  assign _00909_ = w_enq_i & ~(_18408_);
  assign _18409_ = _18390_ | _17487_;
  assign _00910_ = w_enq_i & ~(_18409_);
  assign _18410_ = _18390_ | _17489_;
  assign _00911_ = w_enq_i & ~(_18410_);
  assign _18411_ = _18390_ | _17492_;
  assign _00912_ = w_enq_i & ~(_18411_);
  assign _18412_ = _18390_ | _17494_;
  assign _00913_ = w_enq_i & ~(_18412_);
  assign _18413_ = _18390_ | _17496_;
  assign _00914_ = w_enq_i & ~(_18413_);
  assign _18414_ = _18390_ | _17498_;
  assign _00915_ = w_enq_i & ~(_18414_);
  assign _18415_ = _18390_ | _17502_;
  assign _00916_ = w_enq_i & ~(_18415_);
  assign _18416_ = _18390_ | _17504_;
  assign _00917_ = w_enq_i & ~(_18416_);
  assign _18417_ = _18390_ | _17506_;
  assign _00919_ = w_enq_i & ~(_18417_);
  assign _18418_ = _18390_ | _17508_;
  assign _00920_ = w_enq_i & ~(_18418_);
  assign _18419_ = _18390_ | _17511_;
  assign _00921_ = w_enq_i & ~(_18419_);
  assign _18420_ = _18390_ | _17513_;
  assign _00922_ = w_enq_i & ~(_18420_);
  assign _18421_ = _18390_ | _17515_;
  assign _00923_ = w_enq_i & ~(_18421_);
  assign _18422_ = _18390_ | _17517_;
  assign _00924_ = w_enq_i & ~(_18422_);
  assign _18423_ = _18289_ | _17621_;
  assign _18424_ = _18423_ | _17438_;
  assign _18425_ = _18424_ | _17437_;
  assign _00925_ = w_enq_i & ~(_18425_);
  assign _18426_ = _18424_ | _17444_;
  assign _00926_ = w_enq_i & ~(_18426_);
  assign _18427_ = _18424_ | _17447_;
  assign _00927_ = w_enq_i & ~(_18427_);
  assign _18428_ = _18424_ | _17450_;
  assign _00928_ = w_enq_i & ~(_18428_);
  assign _18429_ = _18424_ | _17454_;
  assign _00931_ = w_enq_i & ~(_18429_);
  assign _18430_ = _18424_ | _17456_;
  assign _00932_ = w_enq_i & ~(_18430_);
  assign _18431_ = _18424_ | _17458_;
  assign _00933_ = w_enq_i & ~(_18431_);
  assign _18432_ = _18424_ | _17460_;
  assign _00934_ = w_enq_i & ~(_18432_);
  assign _18433_ = _18424_ | _17464_;
  assign _00935_ = w_enq_i & ~(_18433_);
  assign _18434_ = _18424_ | _17466_;
  assign _00936_ = w_enq_i & ~(_18434_);
  assign _18435_ = _18424_ | _17468_;
  assign _00937_ = w_enq_i & ~(_18435_);
  assign _18436_ = _18424_ | _17470_;
  assign _00938_ = w_enq_i & ~(_18436_);
  assign _18437_ = _18424_ | _17473_;
  assign _00939_ = w_enq_i & ~(_18437_);
  assign _18438_ = _18424_ | _17475_;
  assign _00940_ = w_enq_i & ~(_18438_);
  assign _18439_ = _18424_ | _17477_;
  assign _00942_ = w_enq_i & ~(_18439_);
  assign _18440_ = _18424_ | _17479_;
  assign _00943_ = w_enq_i & ~(_18440_);
  assign _18441_ = _18424_ | _17483_;
  assign _00944_ = w_enq_i & ~(_18441_);
  assign _18442_ = _18424_ | _17485_;
  assign _00945_ = w_enq_i & ~(_18442_);
  assign _18443_ = _18424_ | _17487_;
  assign _00946_ = w_enq_i & ~(_18443_);
  assign _18444_ = _18424_ | _17489_;
  assign _00947_ = w_enq_i & ~(_18444_);
  assign _18445_ = _18424_ | _17492_;
  assign _00948_ = w_enq_i & ~(_18445_);
  assign _18446_ = _18424_ | _17494_;
  assign _00949_ = w_enq_i & ~(_18446_);
  assign _18447_ = _18424_ | _17496_;
  assign _00950_ = w_enq_i & ~(_18447_);
  assign _18448_ = _18424_ | _17498_;
  assign _00951_ = w_enq_i & ~(_18448_);
  assign _18449_ = _18424_ | _17502_;
  assign _00953_ = w_enq_i & ~(_18449_);
  assign _18450_ = _18424_ | _17504_;
  assign _00954_ = w_enq_i & ~(_18450_);
  assign _18451_ = _18424_ | _17506_;
  assign _00955_ = w_enq_i & ~(_18451_);
  assign _18452_ = _18424_ | _17508_;
  assign _00956_ = w_enq_i & ~(_18452_);
  assign _18453_ = _18424_ | _17511_;
  assign _00957_ = w_enq_i & ~(_18453_);
  assign _18454_ = _18424_ | _17513_;
  assign _00958_ = w_enq_i & ~(_18454_);
  assign _18455_ = _18424_ | _17515_;
  assign _00959_ = w_enq_i & ~(_18455_);
  assign _18456_ = _18424_ | _17517_;
  assign _00960_ = w_enq_i & ~(_18456_);
  assign _18457_ = _18423_ | _17519_;
  assign _18458_ = _18457_ | _17437_;
  assign _00961_ = w_enq_i & ~(_18458_);
  assign _18459_ = _18457_ | _17444_;
  assign _00962_ = w_enq_i & ~(_18459_);
  assign _18460_ = _18457_ | _17447_;
  assign _00964_ = w_enq_i & ~(_18460_);
  assign _18461_ = _18457_ | _17450_;
  assign _00965_ = w_enq_i & ~(_18461_);
  assign _18462_ = _18457_ | _17454_;
  assign _00966_ = w_enq_i & ~(_18462_);
  assign _18463_ = _18457_ | _17456_;
  assign _00967_ = w_enq_i & ~(_18463_);
  assign _18464_ = _18457_ | _17458_;
  assign _00968_ = w_enq_i & ~(_18464_);
  assign _18465_ = _18457_ | _17460_;
  assign _00969_ = w_enq_i & ~(_18465_);
  assign _18466_ = _18457_ | _17464_;
  assign _00970_ = w_enq_i & ~(_18466_);
  assign _18467_ = _18457_ | _17466_;
  assign _00971_ = w_enq_i & ~(_18467_);
  assign _18468_ = _18457_ | _17468_;
  assign _00972_ = w_enq_i & ~(_18468_);
  assign _18469_ = _18457_ | _17470_;
  assign _00973_ = w_enq_i & ~(_18469_);
  assign _18470_ = _18457_ | _17473_;
  assign _00975_ = w_enq_i & ~(_18470_);
  assign _18471_ = _18457_ | _17475_;
  assign _00976_ = w_enq_i & ~(_18471_);
  assign _18472_ = _18457_ | _17477_;
  assign _00977_ = w_enq_i & ~(_18472_);
  assign _18473_ = _18457_ | _17479_;
  assign _00978_ = w_enq_i & ~(_18473_);
  assign _18474_ = _18457_ | _17483_;
  assign _00979_ = w_enq_i & ~(_18474_);
  assign _18475_ = _18457_ | _17485_;
  assign _00980_ = w_enq_i & ~(_18475_);
  assign _18476_ = _18457_ | _17487_;
  assign _00981_ = w_enq_i & ~(_18476_);
  assign _18477_ = _18457_ | _17489_;
  assign _00982_ = w_enq_i & ~(_18477_);
  assign _18478_ = _18457_ | _17492_;
  assign _00983_ = w_enq_i & ~(_18478_);
  assign _18479_ = _18457_ | _17494_;
  assign _00984_ = w_enq_i & ~(_18479_);
  assign _18480_ = _18457_ | _17496_;
  assign _00986_ = w_enq_i & ~(_18480_);
  assign _18481_ = _18457_ | _17498_;
  assign _00987_ = w_enq_i & ~(_18481_);
  assign _18482_ = _18457_ | _17502_;
  assign _00988_ = w_enq_i & ~(_18482_);
  assign _18483_ = _18457_ | _17504_;
  assign _00989_ = w_enq_i & ~(_18483_);
  assign _18484_ = _18457_ | _17506_;
  assign _00990_ = w_enq_i & ~(_18484_);
  assign _18485_ = _18457_ | _17508_;
  assign _00991_ = w_enq_i & ~(_18485_);
  assign _18486_ = _18457_ | _17511_;
  assign _00992_ = w_enq_i & ~(_18486_);
  assign _18487_ = _18457_ | _17513_;
  assign _00993_ = w_enq_i & ~(_18487_);
  assign _18488_ = _18457_ | _17515_;
  assign _00994_ = w_enq_i & ~(_18488_);
  assign _18489_ = _18457_ | _17517_;
  assign _00995_ = w_enq_i & ~(_18489_);
  assign _18490_ = _18423_ | _17553_;
  assign _18491_ = _18490_ | _17437_;
  assign _00997_ = w_enq_i & ~(_18491_);
  assign _18492_ = _18490_ | _17444_;
  assign _00998_ = w_enq_i & ~(_18492_);
  assign _18493_ = _18490_ | _17447_;
  assign _00999_ = w_enq_i & ~(_18493_);
  assign _18494_ = _18490_ | _17450_;
  assign _01000_ = w_enq_i & ~(_18494_);
  assign _18495_ = _18490_ | _17454_;
  assign _01001_ = w_enq_i & ~(_18495_);
  assign _18496_ = _18490_ | _17456_;
  assign _01002_ = w_enq_i & ~(_18496_);
  assign _18497_ = _18490_ | _17458_;
  assign _01003_ = w_enq_i & ~(_18497_);
  assign _18498_ = _18490_ | _17460_;
  assign _01004_ = w_enq_i & ~(_18498_);
  assign _18499_ = _18490_ | _17464_;
  assign _01005_ = w_enq_i & ~(_18499_);
  assign _18500_ = _18490_ | _17466_;
  assign _01006_ = w_enq_i & ~(_18500_);
  assign _18501_ = _18490_ | _17468_;
  assign _01008_ = w_enq_i & ~(_18501_);
  assign _18502_ = _18490_ | _17470_;
  assign _01009_ = w_enq_i & ~(_18502_);
  assign _18503_ = _18490_ | _17473_;
  assign _01010_ = w_enq_i & ~(_18503_);
  assign _18504_ = _18490_ | _17475_;
  assign _01011_ = w_enq_i & ~(_18504_);
  assign _18505_ = _18490_ | _17477_;
  assign _01012_ = w_enq_i & ~(_18505_);
  assign _18506_ = _18490_ | _17479_;
  assign _01013_ = w_enq_i & ~(_18506_);
  assign _18507_ = _18490_ | _17483_;
  assign _01014_ = w_enq_i & ~(_18507_);
  assign _18508_ = _18490_ | _17485_;
  assign _01015_ = w_enq_i & ~(_18508_);
  assign _18509_ = _18490_ | _17487_;
  assign _01016_ = w_enq_i & ~(_18509_);
  assign _18510_ = _18490_ | _17489_;
  assign _01017_ = w_enq_i & ~(_18510_);
  assign _18511_ = _18490_ | _17492_;
  assign _01019_ = w_enq_i & ~(_18511_);
  assign _18512_ = _18490_ | _17494_;
  assign _01020_ = w_enq_i & ~(_18512_);
  assign _18513_ = _18490_ | _17496_;
  assign _01021_ = w_enq_i & ~(_18513_);
  assign _18514_ = _18490_ | _17498_;
  assign _01022_ = w_enq_i & ~(_18514_);
  assign _18515_ = _18490_ | _17502_;
  assign _01023_ = w_enq_i & ~(_18515_);
  assign _18516_ = _18490_ | _17504_;
  assign _01024_ = w_enq_i & ~(_18516_);
  assign _18517_ = _18490_ | _17506_;
  assign _01025_ = w_enq_i & ~(_18517_);
  assign _18518_ = _18490_ | _17508_;
  assign _01026_ = w_enq_i & ~(_18518_);
  assign _18519_ = _18490_ | _17511_;
  assign _01027_ = w_enq_i & ~(_18519_);
  assign _18520_ = _18490_ | _17513_;
  assign _01028_ = w_enq_i & ~(_18520_);
  assign _18521_ = _18490_ | _17515_;
  assign _01030_ = w_enq_i & ~(_18521_);
  assign _18522_ = _18490_ | _17517_;
  assign _01031_ = w_enq_i & ~(_18522_);
  assign _18523_ = _18423_ | _17587_;
  assign _18524_ = _18523_ | _17437_;
  assign _01032_ = w_enq_i & ~(_18524_);
  assign _18525_ = _18523_ | _17444_;
  assign _01033_ = w_enq_i & ~(_18525_);
  assign _18526_ = _18523_ | _17447_;
  assign _01034_ = w_enq_i & ~(_18526_);
  assign _18527_ = _18523_ | _17450_;
  assign _01035_ = w_enq_i & ~(_18527_);
  assign _18528_ = _18523_ | _17454_;
  assign _01036_ = w_enq_i & ~(_18528_);
  assign _18529_ = _18523_ | _17456_;
  assign _01037_ = w_enq_i & ~(_18529_);
  assign _18530_ = _18523_ | _17458_;
  assign _01038_ = w_enq_i & ~(_18530_);
  assign _18531_ = _18523_ | _17460_;
  assign _01039_ = w_enq_i & ~(_18531_);
  assign _18532_ = _18523_ | _17464_;
  assign _00019_ = w_enq_i & ~(_18532_);
  assign _18533_ = _18523_ | _17466_;
  assign _00020_ = w_enq_i & ~(_18533_);
  assign _18534_ = _18523_ | _17468_;
  assign _00021_ = w_enq_i & ~(_18534_);
  assign _18535_ = _18523_ | _17470_;
  assign _00022_ = w_enq_i & ~(_18535_);
  assign _18536_ = _18523_ | _17473_;
  assign _00023_ = w_enq_i & ~(_18536_);
  assign _18537_ = _18523_ | _17475_;
  assign _00024_ = w_enq_i & ~(_18537_);
  assign _18538_ = _18523_ | _17477_;
  assign _00025_ = w_enq_i & ~(_18538_);
  assign _18539_ = _18523_ | _17479_;
  assign _00026_ = w_enq_i & ~(_18539_);
  assign _18540_ = _18523_ | _17483_;
  assign _00027_ = w_enq_i & ~(_18540_);
  assign _18541_ = _18523_ | _17485_;
  assign _00028_ = w_enq_i & ~(_18541_);
  assign _18542_ = _18523_ | _17487_;
  assign _00030_ = w_enq_i & ~(_18542_);
  assign _18543_ = _18523_ | _17489_;
  assign _00031_ = w_enq_i & ~(_18543_);
  assign _18544_ = _18523_ | _17492_;
  assign _00032_ = w_enq_i & ~(_18544_);
  assign _18545_ = _18523_ | _17494_;
  assign _00033_ = w_enq_i & ~(_18545_);
  assign _18546_ = _18523_ | _17496_;
  assign _00034_ = w_enq_i & ~(_18546_);
  assign _18547_ = _18523_ | _17498_;
  assign _00035_ = w_enq_i & ~(_18547_);
  assign _18548_ = _18523_ | _17502_;
  assign _00036_ = w_enq_i & ~(_18548_);
  assign _18549_ = _18523_ | _17504_;
  assign _00037_ = w_enq_i & ~(_18549_);
  assign _18550_ = _18523_ | _17506_;
  assign _00038_ = w_enq_i & ~(_18550_);
  assign _18551_ = _18523_ | _17508_;
  assign _00039_ = w_enq_i & ~(_18551_);
  assign _18552_ = _18523_ | _17511_;
  assign _00041_ = w_enq_i & ~(_18552_);
  assign _18553_ = _18523_ | _17513_;
  assign _00042_ = w_enq_i & ~(_18553_);
  assign _18554_ = _18523_ | _17515_;
  assign _00043_ = w_enq_i & ~(_18554_);
  assign _18555_ = _18523_ | _17517_;
  assign _00044_ = w_enq_i & ~(_18555_);
  assign \bapg_wr.w_ptr_p2 [1] = \bapg_wr.w_ptr_p1_r [1] ^ \bapg_wr.w_ptr_p1_r [0];
  assign _18556_ = \bapg_wr.w_ptr_p1_r [1] & \bapg_wr.w_ptr_p1_r [0];
  assign \bapg_wr.w_ptr_p2 [2] = _18556_ ^ \bapg_wr.w_ptr_p1_r [2];
  assign _18557_ = _18556_ & \bapg_wr.w_ptr_p1_r [2];
  assign \bapg_wr.w_ptr_p2 [3] = _18557_ ^ \bapg_wr.w_ptr_p1_r [3];
  assign _18558_ = ~(\bapg_wr.w_ptr_p1_r [3] & \bapg_wr.w_ptr_p1_r [2]);
  assign _18559_ = _18556_ & ~(_18558_);
  assign \bapg_wr.w_ptr_p2 [4] = _18559_ ^ \bapg_wr.w_ptr_p1_r [4];
  assign _18560_ = _18559_ & \bapg_wr.w_ptr_p1_r [4];
  assign \bapg_wr.w_ptr_p2 [5] = _18560_ ^ \bapg_wr.w_ptr_p1_r [5];
  assign _18561_ = ~(\bapg_wr.w_ptr_p1_r [5] & \bapg_wr.w_ptr_p1_r [4]);
  assign _18562_ = _18559_ & ~(_18561_);
  assign \bapg_wr.w_ptr_p2 [6] = _18562_ ^ \bapg_wr.w_ptr_p1_r [6];
  assign _18563_ = _18562_ & \bapg_wr.w_ptr_p1_r [6];
  assign \bapg_wr.w_ptr_p2 [7] = _18563_ ^ \bapg_wr.w_ptr_p1_r [7];
  assign _18564_ = ~(\bapg_wr.w_ptr_p1_r [7] & \bapg_wr.w_ptr_p1_r [6]);
  assign _18565_ = _18564_ | _18561_;
  assign _18566_ = _18559_ & ~(_18565_);
  assign \bapg_wr.w_ptr_p2 [8] = _18566_ ^ \bapg_wr.w_ptr_p1_r [8];
  assign _18567_ = _18566_ & \bapg_wr.w_ptr_p1_r [8];
  assign \bapg_wr.w_ptr_p2 [9] = _18567_ ^ \bapg_wr.w_ptr_p1_r [9];
  assign _18568_ = ~(\bapg_wr.w_ptr_p1_r [9] & \bapg_wr.w_ptr_p1_r [8]);
  assign _18569_ = _18566_ & ~(_18568_);
  assign \bapg_wr.w_ptr_p2 [10] = _18569_ ^ \bapg_wr.w_ptr_p1_r [10];
  assign \bapg_rd.w_ptr_p2 [1] = \bapg_rd.w_ptr_p1_r [1] ^ \bapg_rd.w_ptr_p1_r [0];
  assign _18570_ = \bapg_rd.w_ptr_p1_r [1] & \bapg_rd.w_ptr_p1_r [0];
  assign \bapg_rd.w_ptr_p2 [2] = _18570_ ^ \bapg_rd.w_ptr_p1_r [2];
  assign _18571_ = _18570_ & \bapg_rd.w_ptr_p1_r [2];
  assign \bapg_rd.w_ptr_p2 [3] = _18571_ ^ \bapg_rd.w_ptr_p1_r [3];
  assign _18572_ = ~(\bapg_rd.w_ptr_p1_r [3] & \bapg_rd.w_ptr_p1_r [2]);
  assign _18573_ = _18570_ & ~(_18572_);
  assign \bapg_rd.w_ptr_p2 [4] = _18573_ ^ \bapg_rd.w_ptr_p1_r [4];
  assign _18574_ = _18573_ & \bapg_rd.w_ptr_p1_r [4];
  assign \bapg_rd.w_ptr_p2 [5] = _18574_ ^ \bapg_rd.w_ptr_p1_r [5];
  assign _18575_ = ~(\bapg_rd.w_ptr_p1_r [5] & \bapg_rd.w_ptr_p1_r [4]);
  assign _18576_ = _18573_ & ~(_18575_);
  assign \bapg_rd.w_ptr_p2 [6] = _18576_ ^ \bapg_rd.w_ptr_p1_r [6];
  assign _18577_ = _18576_ & \bapg_rd.w_ptr_p1_r [6];
  assign \bapg_rd.w_ptr_p2 [7] = _18577_ ^ \bapg_rd.w_ptr_p1_r [7];
  assign _18578_ = ~(\bapg_rd.w_ptr_p1_r [7] & \bapg_rd.w_ptr_p1_r [6]);
  assign _18579_ = _18578_ | _18575_;
  assign _18580_ = _18573_ & ~(_18579_);
  assign \bapg_rd.w_ptr_p2 [8] = _18580_ ^ \bapg_rd.w_ptr_p1_r [8];
  assign _18581_ = _18580_ & \bapg_rd.w_ptr_p1_r [8];
  assign \bapg_rd.w_ptr_p2 [9] = _18581_ ^ \bapg_rd.w_ptr_p1_r [9];
  assign _18582_ = ~(\bapg_rd.w_ptr_p1_r [9] & \bapg_rd.w_ptr_p1_r [8]);
  assign _18583_ = _18580_ & ~(_18582_);
  assign \bapg_rd.w_ptr_p2 [10] = _18583_ ^ \bapg_rd.w_ptr_p1_r [10];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00473_) \MSYNC_1r1w.synth.nz.mem[489] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00462_) \MSYNC_1r1w.synth.nz.mem[479] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00540_) \MSYNC_1r1w.synth.nz.mem[549] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00440_) \MSYNC_1r1w.synth.nz.mem[459] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00451_) \MSYNC_1r1w.synth.nz.mem[469] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00862_) \MSYNC_1r1w.synth.nz.mem[839] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00851_) \MSYNC_1r1w.synth.nz.mem[829] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00529_) \MSYNC_1r1w.synth.nz.mem[539] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00429_) \MSYNC_1r1w.synth.nz.mem[449] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00518_) \MSYNC_1r1w.synth.nz.mem[529] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00418_) \MSYNC_1r1w.synth.nz.mem[439] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00662_) \MSYNC_1r1w.synth.nz.mem[659] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00629_) \MSYNC_1r1w.synth.nz.mem[629] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00618_) \MSYNC_1r1w.synth.nz.mem[619] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00607_) \MSYNC_1r1w.synth.nz.mem[609] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00673_) \MSYNC_1r1w.synth.nz.mem[669] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00595_) \MSYNC_1r1w.synth.nz.mem[599] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01017_) \MSYNC_1r1w.synth.nz.mem[979] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00584_) \MSYNC_1r1w.synth.nz.mem[589] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00573_) \MSYNC_1r1w.synth.nz.mem[579] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00806_) \MSYNC_1r1w.synth.nz.mem[789] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00884_) \MSYNC_1r1w.synth.nz.mem[859] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00840_) \MSYNC_1r1w.synth.nz.mem[819] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00829_) \MSYNC_1r1w.synth.nz.mem[809] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01006_) \MSYNC_1r1w.synth.nz.mem[969] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00895_) \MSYNC_1r1w.synth.nz.mem[869] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00951_) \MSYNC_1r1w.synth.nz.mem[919] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00196_) \MSYNC_1r1w.synth.nz.mem[239] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00917_) \MSYNC_1r1w.synth.nz.mem[889] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00817_) \MSYNC_1r1w.synth.nz.mem[799] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00562_) \MSYNC_1r1w.synth.nz.mem[569] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00651_) \MSYNC_1r1w.synth.nz.mem[649] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00551_) \MSYNC_1r1w.synth.nz.mem[559] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00407_) \MSYNC_1r1w.synth.nz.mem[429] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00396_) \MSYNC_1r1w.synth.nz.mem[419] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00507_) \MSYNC_1r1w.synth.nz.mem[519] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00906_) \MSYNC_1r1w.synth.nz.mem[879] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00873_) \MSYNC_1r1w.synth.nz.mem[849] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00640_) \MSYNC_1r1w.synth.nz.mem[639] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00995_) \MSYNC_1r1w.synth.nz.mem[959] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00962_) \MSYNC_1r1w.synth.nz.mem[929] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00984_) \MSYNC_1r1w.synth.nz.mem[949] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00973_) \MSYNC_1r1w.synth.nz.mem[939] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01039_) \MSYNC_1r1w.synth.nz.mem[999] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00373_) \MSYNC_1r1w.synth.nz.mem[399] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00940_) \MSYNC_1r1w.synth.nz.mem[909] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00385_) \MSYNC_1r1w.synth.nz.mem[409] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00928_) \MSYNC_1r1w.synth.nz.mem[899] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01028_) \MSYNC_1r1w.synth.nz.mem[989] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00028_) \MSYNC_1r1w.synth.nz.mem[1009] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00362_) \MSYNC_1r1w.synth.nz.mem[389] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00351_) \MSYNC_1r1w.synth.nz.mem[379] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00340_) \MSYNC_1r1w.synth.nz.mem[369] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00329_) \MSYNC_1r1w.synth.nz.mem[359] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00318_) \MSYNC_1r1w.synth.nz.mem[349] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00307_) \MSYNC_1r1w.synth.nz.mem[339] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00296_) \MSYNC_1r1w.synth.nz.mem[329] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00762_) \MSYNC_1r1w.synth.nz.mem[749] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00285_) \MSYNC_1r1w.synth.nz.mem[319] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00773_) \MSYNC_1r1w.synth.nz.mem[759] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00274_) \MSYNC_1r1w.synth.nz.mem[309] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00496_) \MSYNC_1r1w.synth.nz.mem[509] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00484_) \MSYNC_1r1w.synth.nz.mem[499] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00751_) \MSYNC_1r1w.synth.nz.mem[739] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00740_) \MSYNC_1r1w.synth.nz.mem[729] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00729_) \MSYNC_1r1w.synth.nz.mem[719] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00718_) \MSYNC_1r1w.synth.nz.mem[709] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00706_) \MSYNC_1r1w.synth.nz.mem[699] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00695_) \MSYNC_1r1w.synth.nz.mem[689] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00684_) \MSYNC_1r1w.synth.nz.mem[679] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00795_) \MSYNC_1r1w.synth.nz.mem[779] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00784_) \MSYNC_1r1w.synth.nz.mem[769] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00251_) \MSYNC_1r1w.synth.nz.mem[289] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00240_) \MSYNC_1r1w.synth.nz.mem[279] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00152_) \MSYNC_1r1w.synth.nz.mem[19] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00229_) \MSYNC_1r1w.synth.nz.mem[269] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00218_) \MSYNC_1r1w.synth.nz.mem[259] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00207_) \MSYNC_1r1w.synth.nz.mem[249] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00818_) \MSYNC_1r1w.synth.nz.mem[79] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00262_) \MSYNC_1r1w.synth.nz.mem[299] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00185_) \MSYNC_1r1w.synth.nz.mem[229] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00174_) \MSYNC_1r1w.synth.nz.mem[219] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00163_) \MSYNC_1r1w.synth.nz.mem[209] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00596_) \MSYNC_1r1w.synth.nz.mem[59] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00263_) \MSYNC_1r1w.synth.nz.mem[29] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00151_) \MSYNC_1r1w.synth.nz.mem[199] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00374_) \MSYNC_1r1w.synth.nz.mem[39] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00140_) \MSYNC_1r1w.synth.nz.mem[189] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00707_) \MSYNC_1r1w.synth.nz.mem[69] [15] <= w_data_i[15];
  reg \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[1] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[1]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[1]  <= _00000_;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [1] = \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[1] ;
  reg \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[2] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[2]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[2]  <= _00001_;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [2] = \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[2] ;
  reg \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[3] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[3]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[3]  <= _00002_;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [3] = \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[3] ;
  reg \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[4] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[4]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[4]  <= _00003_;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [4] = \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[4] ;
  reg \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[5] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[5]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[5]  <= _00004_;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [5] = \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[5] ;
  reg \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[6] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[6]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[6]  <= _00005_;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [6] = \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[6] ;
  reg \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[7] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[7]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[7]  <= _00006_;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7] = \bapg_wr.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[7] ;
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [0] <= \bapg_wr.w_ptr_p1_r [1];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [1] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [1];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [2] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [2];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [3] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [3];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [4] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [4];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [5] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [5];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [6] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [6];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [7] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [0] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [0];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [1] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [1];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [2] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [2];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [3] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [3];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [4] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [4];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [5] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [5];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [6] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [6];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [7] <= \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [7];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= _00007_;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= _00008_;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [2] <= 1'h0;
    else if (w_enq_i) \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [2] <= \bapg_wr.w_ptr_p1_r [10];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0] <= \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1] <= \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [2] <= \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [2];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] <= \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] <= \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1];
  always @(posedge r_clk_i)
    \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [2] <= \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [2];
  reg \bapg_wr.w_ptr_r_reg[0] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[0]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[0]  <= \bapg_wr.w_ptr_p1_r [0];
  assign \bapg_wr.w_ptr_r [0] = \bapg_wr.w_ptr_r_reg[0] ;
  reg \bapg_wr.w_ptr_r_reg[1] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[1]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[1]  <= \bapg_wr.w_ptr_p1_r [1];
  assign \bapg_wr.w_ptr_r [1] = \bapg_wr.w_ptr_r_reg[1] ;
  reg \bapg_wr.w_ptr_r_reg[2] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[2]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[2]  <= \bapg_wr.w_ptr_p1_r [2];
  assign \bapg_wr.w_ptr_r [2] = \bapg_wr.w_ptr_r_reg[2] ;
  reg \bapg_wr.w_ptr_r_reg[3] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[3]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[3]  <= \bapg_wr.w_ptr_p1_r [3];
  assign \bapg_wr.w_ptr_r [3] = \bapg_wr.w_ptr_r_reg[3] ;
  reg \bapg_wr.w_ptr_r_reg[4] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[4]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[4]  <= \bapg_wr.w_ptr_p1_r [4];
  assign \bapg_wr.w_ptr_r [4] = \bapg_wr.w_ptr_r_reg[4] ;
  reg \bapg_wr.w_ptr_r_reg[5] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[5]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[5]  <= \bapg_wr.w_ptr_p1_r [5];
  assign \bapg_wr.w_ptr_r [5] = \bapg_wr.w_ptr_r_reg[5] ;
  reg \bapg_wr.w_ptr_r_reg[6] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[6]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[6]  <= \bapg_wr.w_ptr_p1_r [6];
  assign \bapg_wr.w_ptr_r [6] = \bapg_wr.w_ptr_r_reg[6] ;
  reg \bapg_wr.w_ptr_r_reg[7] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[7]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[7]  <= \bapg_wr.w_ptr_p1_r [7];
  assign \bapg_wr.w_ptr_r [7] = \bapg_wr.w_ptr_r_reg[7] ;
  reg \bapg_wr.w_ptr_r_reg[8] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[8]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[8]  <= \bapg_wr.w_ptr_p1_r [8];
  assign \bapg_wr.w_ptr_r [8] = \bapg_wr.w_ptr_r_reg[8] ;
  reg \bapg_wr.w_ptr_r_reg[9] ;
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_r_reg[9]  <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_r_reg[9]  <= \bapg_wr.w_ptr_p1_r [9];
  assign \bapg_wr.w_ptr_r [9] = \bapg_wr.w_ptr_r_reg[9] ;
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00074_) \MSYNC_1r1w.synth.nz.mem[129] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [0] <= 1'h1;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [0] <= \bapg_wr.w_ptr_p2 [0];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [1] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [1] <= \bapg_wr.w_ptr_p2 [1];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [2] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [2] <= \bapg_wr.w_ptr_p2 [2];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [3] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [3] <= \bapg_wr.w_ptr_p2 [3];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [4] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [4] <= \bapg_wr.w_ptr_p2 [4];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [5] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [5] <= \bapg_wr.w_ptr_p2 [5];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [6] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [6] <= \bapg_wr.w_ptr_p2 [6];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [7] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [7] <= \bapg_wr.w_ptr_p2 [7];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [8] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [8] <= \bapg_wr.w_ptr_p2 [8];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [9] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [9] <= \bapg_wr.w_ptr_p2 [9];
  always @(posedge w_clk_i)
    if (w_reset_i) \bapg_wr.w_ptr_p1_r [10] <= 1'h0;
    else if (w_enq_i) \bapg_wr.w_ptr_p1_r [10] <= \bapg_wr.w_ptr_p2 [10];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00063_) \MSYNC_1r1w.synth.nz.mem[119] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00129_) \MSYNC_1r1w.synth.nz.mem[179] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00485_) \MSYNC_1r1w.synth.nz.mem[49] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00118_) \MSYNC_1r1w.synth.nz.mem[169] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00107_) \MSYNC_1r1w.synth.nz.mem[159] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00096_) \MSYNC_1r1w.synth.nz.mem[149] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00085_) \MSYNC_1r1w.synth.nz.mem[139] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00045_) \MSYNC_1r1w.synth.nz.mem[102] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00044_) \MSYNC_1r1w.synth.nz.mem[1023] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00039_) \MSYNC_1r1w.synth.nz.mem[1019] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00052_) \MSYNC_1r1w.synth.nz.mem[109] [15] <= w_data_i[15];
  reg \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[1] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[1]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[1]  <= _00009_;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [1] = \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[1] ;
  reg \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[2] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[2]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[2]  <= _00010_;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [2] = \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[2] ;
  reg \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[3] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[3]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[3]  <= _00011_;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [3] = \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[3] ;
  reg \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[4] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[4]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[4]  <= _00012_;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [4] = \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[4] ;
  reg \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[5] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[5]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[5]  <= _00013_;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [5] = \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[5] ;
  reg \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[6] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[6]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[6]  <= _00014_;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [6] = \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[6] ;
  reg \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[7] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[7]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[7]  <= _00015_;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7] = \bapg_rd.ptr_sync.sync.p.maxb_reg[0].blss.bsg_SYNC_LNCH_r[7] ;
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [0] <= \bapg_rd.w_ptr_p1_r [1];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [1] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [1];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [2] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [2];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [3] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [3];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [4] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [4];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [5] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [5];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [6] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [6];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [7] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [0] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [0];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [1] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [1];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [2] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [2];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [3] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [3];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [4] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [4];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [5] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [5];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [6] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [6];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r [7] <= \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_1_r [7];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0] <= _00016_;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1] <= _00017_;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [2] <= 1'h0;
    else if (r_deq_i) \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [2] <= \bapg_rd.w_ptr_p1_r [10];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0] <= \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [0];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1] <= \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [1];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [2] <= \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r [2];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [0] <= \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [0];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [1] <= \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [1];
  always @(posedge w_clk_i)
    \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r [2] <= \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_1_r [2];
  reg \bapg_rd.w_ptr_r_reg[0] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[0]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[0]  <= \bapg_rd.w_ptr_p1_r [0];
  assign \bapg_rd.w_ptr_r [0] = \bapg_rd.w_ptr_r_reg[0] ;
  reg \bapg_rd.w_ptr_r_reg[1] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[1]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[1]  <= \bapg_rd.w_ptr_p1_r [1];
  assign \bapg_rd.w_ptr_r [1] = \bapg_rd.w_ptr_r_reg[1] ;
  reg \bapg_rd.w_ptr_r_reg[2] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[2]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[2]  <= \bapg_rd.w_ptr_p1_r [2];
  assign \bapg_rd.w_ptr_r [2] = \bapg_rd.w_ptr_r_reg[2] ;
  reg \bapg_rd.w_ptr_r_reg[3] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[3]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[3]  <= \bapg_rd.w_ptr_p1_r [3];
  assign \bapg_rd.w_ptr_r [3] = \bapg_rd.w_ptr_r_reg[3] ;
  reg \bapg_rd.w_ptr_r_reg[4] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[4]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[4]  <= \bapg_rd.w_ptr_p1_r [4];
  assign \bapg_rd.w_ptr_r [4] = \bapg_rd.w_ptr_r_reg[4] ;
  reg \bapg_rd.w_ptr_r_reg[5] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[5]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[5]  <= \bapg_rd.w_ptr_p1_r [5];
  assign \bapg_rd.w_ptr_r [5] = \bapg_rd.w_ptr_r_reg[5] ;
  reg \bapg_rd.w_ptr_r_reg[6] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[6]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[6]  <= \bapg_rd.w_ptr_p1_r [6];
  assign \bapg_rd.w_ptr_r [6] = \bapg_rd.w_ptr_r_reg[6] ;
  reg \bapg_rd.w_ptr_r_reg[7] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[7]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[7]  <= \bapg_rd.w_ptr_p1_r [7];
  assign \bapg_rd.w_ptr_r [7] = \bapg_rd.w_ptr_r_reg[7] ;
  reg \bapg_rd.w_ptr_r_reg[8] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[8]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[8]  <= \bapg_rd.w_ptr_p1_r [8];
  assign \bapg_rd.w_ptr_r [8] = \bapg_rd.w_ptr_r_reg[8] ;
  reg \bapg_rd.w_ptr_r_reg[9] ;
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_r_reg[9]  <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_r_reg[9]  <= \bapg_rd.w_ptr_p1_r [9];
  assign \bapg_rd.w_ptr_r [9] = \bapg_rd.w_ptr_r_reg[9] ;
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01040_) \MSYNC_1r1w.synth.nz.mem[99] [15] <= w_data_i[15];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [0] <= 1'h1;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [0] <= \bapg_rd.w_ptr_p2 [0];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [1] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [1] <= \bapg_rd.w_ptr_p2 [1];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [2] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [2] <= \bapg_rd.w_ptr_p2 [2];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [3] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [3] <= \bapg_rd.w_ptr_p2 [3];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [4] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [4] <= \bapg_rd.w_ptr_p2 [4];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [5] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [5] <= \bapg_rd.w_ptr_p2 [5];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [6] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [6] <= \bapg_rd.w_ptr_p2 [6];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [7] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [7] <= \bapg_rd.w_ptr_p2 [7];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [8] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [8] <= \bapg_rd.w_ptr_p2 [8];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [9] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [9] <= \bapg_rd.w_ptr_p2 [9];
  always @(posedge r_clk_i)
    if (r_reset_i) \bapg_rd.w_ptr_p1_r [10] <= 1'h0;
    else if (r_deq_i) \bapg_rd.w_ptr_p1_r [10] <= \bapg_rd.w_ptr_p2 [10];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00929_) \MSYNC_1r1w.synth.nz.mem[89] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00046_) \MSYNC_1r1w.synth.nz.mem[103] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00047_) \MSYNC_1r1w.synth.nz.mem[104] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00048_) \MSYNC_1r1w.synth.nz.mem[105] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00049_) \MSYNC_1r1w.synth.nz.mem[106] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00050_) \MSYNC_1r1w.synth.nz.mem[107] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00051_) \MSYNC_1r1w.synth.nz.mem[108] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00053_) \MSYNC_1r1w.synth.nz.mem[10] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00054_) \MSYNC_1r1w.synth.nz.mem[110] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00055_) \MSYNC_1r1w.synth.nz.mem[111] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00056_) \MSYNC_1r1w.synth.nz.mem[112] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00057_) \MSYNC_1r1w.synth.nz.mem[113] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00058_) \MSYNC_1r1w.synth.nz.mem[114] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00059_) \MSYNC_1r1w.synth.nz.mem[115] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00060_) \MSYNC_1r1w.synth.nz.mem[116] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00061_) \MSYNC_1r1w.synth.nz.mem[117] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00062_) \MSYNC_1r1w.synth.nz.mem[118] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00064_) \MSYNC_1r1w.synth.nz.mem[11] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00065_) \MSYNC_1r1w.synth.nz.mem[120] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00066_) \MSYNC_1r1w.synth.nz.mem[121] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00067_) \MSYNC_1r1w.synth.nz.mem[122] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00068_) \MSYNC_1r1w.synth.nz.mem[123] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00069_) \MSYNC_1r1w.synth.nz.mem[124] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00070_) \MSYNC_1r1w.synth.nz.mem[125] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00071_) \MSYNC_1r1w.synth.nz.mem[126] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00072_) \MSYNC_1r1w.synth.nz.mem[127] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00073_) \MSYNC_1r1w.synth.nz.mem[128] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00075_) \MSYNC_1r1w.synth.nz.mem[12] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00076_) \MSYNC_1r1w.synth.nz.mem[130] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00077_) \MSYNC_1r1w.synth.nz.mem[131] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00078_) \MSYNC_1r1w.synth.nz.mem[132] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00079_) \MSYNC_1r1w.synth.nz.mem[133] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00080_) \MSYNC_1r1w.synth.nz.mem[134] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00081_) \MSYNC_1r1w.synth.nz.mem[135] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00082_) \MSYNC_1r1w.synth.nz.mem[136] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00083_) \MSYNC_1r1w.synth.nz.mem[137] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00084_) \MSYNC_1r1w.synth.nz.mem[138] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00086_) \MSYNC_1r1w.synth.nz.mem[13] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00087_) \MSYNC_1r1w.synth.nz.mem[140] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00088_) \MSYNC_1r1w.synth.nz.mem[141] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00089_) \MSYNC_1r1w.synth.nz.mem[142] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00090_) \MSYNC_1r1w.synth.nz.mem[143] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00091_) \MSYNC_1r1w.synth.nz.mem[144] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00092_) \MSYNC_1r1w.synth.nz.mem[145] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00093_) \MSYNC_1r1w.synth.nz.mem[146] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00094_) \MSYNC_1r1w.synth.nz.mem[147] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00095_) \MSYNC_1r1w.synth.nz.mem[148] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00097_) \MSYNC_1r1w.synth.nz.mem[14] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00098_) \MSYNC_1r1w.synth.nz.mem[150] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00099_) \MSYNC_1r1w.synth.nz.mem[151] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00100_) \MSYNC_1r1w.synth.nz.mem[152] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00101_) \MSYNC_1r1w.synth.nz.mem[153] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00102_) \MSYNC_1r1w.synth.nz.mem[154] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00103_) \MSYNC_1r1w.synth.nz.mem[155] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00104_) \MSYNC_1r1w.synth.nz.mem[156] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00105_) \MSYNC_1r1w.synth.nz.mem[157] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00106_) \MSYNC_1r1w.synth.nz.mem[158] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00108_) \MSYNC_1r1w.synth.nz.mem[15] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00109_) \MSYNC_1r1w.synth.nz.mem[160] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00110_) \MSYNC_1r1w.synth.nz.mem[161] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00111_) \MSYNC_1r1w.synth.nz.mem[162] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00112_) \MSYNC_1r1w.synth.nz.mem[163] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00113_) \MSYNC_1r1w.synth.nz.mem[164] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00114_) \MSYNC_1r1w.synth.nz.mem[165] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00115_) \MSYNC_1r1w.synth.nz.mem[166] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00116_) \MSYNC_1r1w.synth.nz.mem[167] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00117_) \MSYNC_1r1w.synth.nz.mem[168] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00119_) \MSYNC_1r1w.synth.nz.mem[16] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00120_) \MSYNC_1r1w.synth.nz.mem[170] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00121_) \MSYNC_1r1w.synth.nz.mem[171] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00122_) \MSYNC_1r1w.synth.nz.mem[172] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00123_) \MSYNC_1r1w.synth.nz.mem[173] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00124_) \MSYNC_1r1w.synth.nz.mem[174] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00125_) \MSYNC_1r1w.synth.nz.mem[175] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00126_) \MSYNC_1r1w.synth.nz.mem[176] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00127_) \MSYNC_1r1w.synth.nz.mem[177] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00128_) \MSYNC_1r1w.synth.nz.mem[178] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00130_) \MSYNC_1r1w.synth.nz.mem[17] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00131_) \MSYNC_1r1w.synth.nz.mem[180] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00132_) \MSYNC_1r1w.synth.nz.mem[181] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00133_) \MSYNC_1r1w.synth.nz.mem[182] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00134_) \MSYNC_1r1w.synth.nz.mem[183] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00135_) \MSYNC_1r1w.synth.nz.mem[184] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00136_) \MSYNC_1r1w.synth.nz.mem[185] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00137_) \MSYNC_1r1w.synth.nz.mem[186] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00138_) \MSYNC_1r1w.synth.nz.mem[187] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00139_) \MSYNC_1r1w.synth.nz.mem[188] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00141_) \MSYNC_1r1w.synth.nz.mem[18] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00142_) \MSYNC_1r1w.synth.nz.mem[190] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00143_) \MSYNC_1r1w.synth.nz.mem[191] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00144_) \MSYNC_1r1w.synth.nz.mem[192] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00145_) \MSYNC_1r1w.synth.nz.mem[193] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00146_) \MSYNC_1r1w.synth.nz.mem[194] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00147_) \MSYNC_1r1w.synth.nz.mem[195] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00148_) \MSYNC_1r1w.synth.nz.mem[196] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00149_) \MSYNC_1r1w.synth.nz.mem[197] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00150_) \MSYNC_1r1w.synth.nz.mem[198] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00153_) \MSYNC_1r1w.synth.nz.mem[1] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00154_) \MSYNC_1r1w.synth.nz.mem[200] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00155_) \MSYNC_1r1w.synth.nz.mem[201] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00156_) \MSYNC_1r1w.synth.nz.mem[202] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00157_) \MSYNC_1r1w.synth.nz.mem[203] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00158_) \MSYNC_1r1w.synth.nz.mem[204] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00159_) \MSYNC_1r1w.synth.nz.mem[205] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00160_) \MSYNC_1r1w.synth.nz.mem[206] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00161_) \MSYNC_1r1w.synth.nz.mem[207] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00162_) \MSYNC_1r1w.synth.nz.mem[208] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00164_) \MSYNC_1r1w.synth.nz.mem[20] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00165_) \MSYNC_1r1w.synth.nz.mem[210] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00166_) \MSYNC_1r1w.synth.nz.mem[211] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00167_) \MSYNC_1r1w.synth.nz.mem[212] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00168_) \MSYNC_1r1w.synth.nz.mem[213] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00169_) \MSYNC_1r1w.synth.nz.mem[214] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00170_) \MSYNC_1r1w.synth.nz.mem[215] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00171_) \MSYNC_1r1w.synth.nz.mem[216] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00172_) \MSYNC_1r1w.synth.nz.mem[217] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00173_) \MSYNC_1r1w.synth.nz.mem[218] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00175_) \MSYNC_1r1w.synth.nz.mem[21] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00176_) \MSYNC_1r1w.synth.nz.mem[220] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00177_) \MSYNC_1r1w.synth.nz.mem[221] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00178_) \MSYNC_1r1w.synth.nz.mem[222] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00179_) \MSYNC_1r1w.synth.nz.mem[223] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00180_) \MSYNC_1r1w.synth.nz.mem[224] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00181_) \MSYNC_1r1w.synth.nz.mem[225] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00182_) \MSYNC_1r1w.synth.nz.mem[226] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00183_) \MSYNC_1r1w.synth.nz.mem[227] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00184_) \MSYNC_1r1w.synth.nz.mem[228] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00186_) \MSYNC_1r1w.synth.nz.mem[22] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00187_) \MSYNC_1r1w.synth.nz.mem[230] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00188_) \MSYNC_1r1w.synth.nz.mem[231] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00189_) \MSYNC_1r1w.synth.nz.mem[232] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00190_) \MSYNC_1r1w.synth.nz.mem[233] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00191_) \MSYNC_1r1w.synth.nz.mem[234] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00192_) \MSYNC_1r1w.synth.nz.mem[235] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00193_) \MSYNC_1r1w.synth.nz.mem[236] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00194_) \MSYNC_1r1w.synth.nz.mem[237] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00195_) \MSYNC_1r1w.synth.nz.mem[238] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00197_) \MSYNC_1r1w.synth.nz.mem[23] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00198_) \MSYNC_1r1w.synth.nz.mem[240] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00199_) \MSYNC_1r1w.synth.nz.mem[241] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00200_) \MSYNC_1r1w.synth.nz.mem[242] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00201_) \MSYNC_1r1w.synth.nz.mem[243] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00202_) \MSYNC_1r1w.synth.nz.mem[244] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00203_) \MSYNC_1r1w.synth.nz.mem[245] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00204_) \MSYNC_1r1w.synth.nz.mem[246] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00205_) \MSYNC_1r1w.synth.nz.mem[247] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00206_) \MSYNC_1r1w.synth.nz.mem[248] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00208_) \MSYNC_1r1w.synth.nz.mem[24] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00209_) \MSYNC_1r1w.synth.nz.mem[250] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00210_) \MSYNC_1r1w.synth.nz.mem[251] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00211_) \MSYNC_1r1w.synth.nz.mem[252] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00212_) \MSYNC_1r1w.synth.nz.mem[253] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00213_) \MSYNC_1r1w.synth.nz.mem[254] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00214_) \MSYNC_1r1w.synth.nz.mem[255] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00215_) \MSYNC_1r1w.synth.nz.mem[256] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00216_) \MSYNC_1r1w.synth.nz.mem[257] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00217_) \MSYNC_1r1w.synth.nz.mem[258] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00219_) \MSYNC_1r1w.synth.nz.mem[25] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00220_) \MSYNC_1r1w.synth.nz.mem[260] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00221_) \MSYNC_1r1w.synth.nz.mem[261] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00222_) \MSYNC_1r1w.synth.nz.mem[262] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00223_) \MSYNC_1r1w.synth.nz.mem[263] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00224_) \MSYNC_1r1w.synth.nz.mem[264] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00225_) \MSYNC_1r1w.synth.nz.mem[265] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00226_) \MSYNC_1r1w.synth.nz.mem[266] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00227_) \MSYNC_1r1w.synth.nz.mem[267] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00228_) \MSYNC_1r1w.synth.nz.mem[268] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00230_) \MSYNC_1r1w.synth.nz.mem[26] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00231_) \MSYNC_1r1w.synth.nz.mem[270] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00232_) \MSYNC_1r1w.synth.nz.mem[271] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00233_) \MSYNC_1r1w.synth.nz.mem[272] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00234_) \MSYNC_1r1w.synth.nz.mem[273] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00235_) \MSYNC_1r1w.synth.nz.mem[274] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00236_) \MSYNC_1r1w.synth.nz.mem[275] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00237_) \MSYNC_1r1w.synth.nz.mem[276] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00238_) \MSYNC_1r1w.synth.nz.mem[277] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00239_) \MSYNC_1r1w.synth.nz.mem[278] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00241_) \MSYNC_1r1w.synth.nz.mem[27] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00242_) \MSYNC_1r1w.synth.nz.mem[280] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00243_) \MSYNC_1r1w.synth.nz.mem[281] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00244_) \MSYNC_1r1w.synth.nz.mem[282] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00245_) \MSYNC_1r1w.synth.nz.mem[283] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00246_) \MSYNC_1r1w.synth.nz.mem[284] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00247_) \MSYNC_1r1w.synth.nz.mem[285] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00248_) \MSYNC_1r1w.synth.nz.mem[286] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00249_) \MSYNC_1r1w.synth.nz.mem[287] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00250_) \MSYNC_1r1w.synth.nz.mem[288] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00252_) \MSYNC_1r1w.synth.nz.mem[28] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00253_) \MSYNC_1r1w.synth.nz.mem[290] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00254_) \MSYNC_1r1w.synth.nz.mem[291] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00255_) \MSYNC_1r1w.synth.nz.mem[292] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00256_) \MSYNC_1r1w.synth.nz.mem[293] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00257_) \MSYNC_1r1w.synth.nz.mem[294] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00258_) \MSYNC_1r1w.synth.nz.mem[295] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00259_) \MSYNC_1r1w.synth.nz.mem[296] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00260_) \MSYNC_1r1w.synth.nz.mem[297] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00261_) \MSYNC_1r1w.synth.nz.mem[298] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00264_) \MSYNC_1r1w.synth.nz.mem[2] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00265_) \MSYNC_1r1w.synth.nz.mem[300] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00266_) \MSYNC_1r1w.synth.nz.mem[301] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00267_) \MSYNC_1r1w.synth.nz.mem[302] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00268_) \MSYNC_1r1w.synth.nz.mem[303] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00269_) \MSYNC_1r1w.synth.nz.mem[304] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00270_) \MSYNC_1r1w.synth.nz.mem[305] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00271_) \MSYNC_1r1w.synth.nz.mem[306] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00272_) \MSYNC_1r1w.synth.nz.mem[307] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00273_) \MSYNC_1r1w.synth.nz.mem[308] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00275_) \MSYNC_1r1w.synth.nz.mem[30] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00276_) \MSYNC_1r1w.synth.nz.mem[310] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00277_) \MSYNC_1r1w.synth.nz.mem[311] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00278_) \MSYNC_1r1w.synth.nz.mem[312] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00279_) \MSYNC_1r1w.synth.nz.mem[313] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00280_) \MSYNC_1r1w.synth.nz.mem[314] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00281_) \MSYNC_1r1w.synth.nz.mem[315] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00282_) \MSYNC_1r1w.synth.nz.mem[316] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00283_) \MSYNC_1r1w.synth.nz.mem[317] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00284_) \MSYNC_1r1w.synth.nz.mem[318] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00286_) \MSYNC_1r1w.synth.nz.mem[31] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00287_) \MSYNC_1r1w.synth.nz.mem[320] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00288_) \MSYNC_1r1w.synth.nz.mem[321] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00289_) \MSYNC_1r1w.synth.nz.mem[322] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00290_) \MSYNC_1r1w.synth.nz.mem[323] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00291_) \MSYNC_1r1w.synth.nz.mem[324] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00292_) \MSYNC_1r1w.synth.nz.mem[325] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00293_) \MSYNC_1r1w.synth.nz.mem[326] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00294_) \MSYNC_1r1w.synth.nz.mem[327] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00295_) \MSYNC_1r1w.synth.nz.mem[328] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00297_) \MSYNC_1r1w.synth.nz.mem[32] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00298_) \MSYNC_1r1w.synth.nz.mem[330] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00299_) \MSYNC_1r1w.synth.nz.mem[331] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00300_) \MSYNC_1r1w.synth.nz.mem[332] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00301_) \MSYNC_1r1w.synth.nz.mem[333] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00302_) \MSYNC_1r1w.synth.nz.mem[334] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00303_) \MSYNC_1r1w.synth.nz.mem[335] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00304_) \MSYNC_1r1w.synth.nz.mem[336] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00305_) \MSYNC_1r1w.synth.nz.mem[337] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00306_) \MSYNC_1r1w.synth.nz.mem[338] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00308_) \MSYNC_1r1w.synth.nz.mem[33] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00309_) \MSYNC_1r1w.synth.nz.mem[340] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00310_) \MSYNC_1r1w.synth.nz.mem[341] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00311_) \MSYNC_1r1w.synth.nz.mem[342] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00312_) \MSYNC_1r1w.synth.nz.mem[343] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00313_) \MSYNC_1r1w.synth.nz.mem[344] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00314_) \MSYNC_1r1w.synth.nz.mem[345] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00315_) \MSYNC_1r1w.synth.nz.mem[346] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00316_) \MSYNC_1r1w.synth.nz.mem[347] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00317_) \MSYNC_1r1w.synth.nz.mem[348] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00319_) \MSYNC_1r1w.synth.nz.mem[34] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00320_) \MSYNC_1r1w.synth.nz.mem[350] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00321_) \MSYNC_1r1w.synth.nz.mem[351] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00322_) \MSYNC_1r1w.synth.nz.mem[352] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00323_) \MSYNC_1r1w.synth.nz.mem[353] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00324_) \MSYNC_1r1w.synth.nz.mem[354] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00325_) \MSYNC_1r1w.synth.nz.mem[355] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00326_) \MSYNC_1r1w.synth.nz.mem[356] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00327_) \MSYNC_1r1w.synth.nz.mem[357] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00328_) \MSYNC_1r1w.synth.nz.mem[358] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00330_) \MSYNC_1r1w.synth.nz.mem[35] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00331_) \MSYNC_1r1w.synth.nz.mem[360] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00332_) \MSYNC_1r1w.synth.nz.mem[361] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00333_) \MSYNC_1r1w.synth.nz.mem[362] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00334_) \MSYNC_1r1w.synth.nz.mem[363] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00335_) \MSYNC_1r1w.synth.nz.mem[364] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00336_) \MSYNC_1r1w.synth.nz.mem[365] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00337_) \MSYNC_1r1w.synth.nz.mem[366] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00338_) \MSYNC_1r1w.synth.nz.mem[367] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00339_) \MSYNC_1r1w.synth.nz.mem[368] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00341_) \MSYNC_1r1w.synth.nz.mem[36] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00342_) \MSYNC_1r1w.synth.nz.mem[370] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00343_) \MSYNC_1r1w.synth.nz.mem[371] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00344_) \MSYNC_1r1w.synth.nz.mem[372] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00345_) \MSYNC_1r1w.synth.nz.mem[373] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00346_) \MSYNC_1r1w.synth.nz.mem[374] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00347_) \MSYNC_1r1w.synth.nz.mem[375] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00348_) \MSYNC_1r1w.synth.nz.mem[376] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00349_) \MSYNC_1r1w.synth.nz.mem[377] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00350_) \MSYNC_1r1w.synth.nz.mem[378] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00352_) \MSYNC_1r1w.synth.nz.mem[37] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00353_) \MSYNC_1r1w.synth.nz.mem[380] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00354_) \MSYNC_1r1w.synth.nz.mem[381] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00355_) \MSYNC_1r1w.synth.nz.mem[382] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00356_) \MSYNC_1r1w.synth.nz.mem[383] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00357_) \MSYNC_1r1w.synth.nz.mem[384] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00358_) \MSYNC_1r1w.synth.nz.mem[385] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00359_) \MSYNC_1r1w.synth.nz.mem[386] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00360_) \MSYNC_1r1w.synth.nz.mem[387] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00361_) \MSYNC_1r1w.synth.nz.mem[388] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00363_) \MSYNC_1r1w.synth.nz.mem[38] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00364_) \MSYNC_1r1w.synth.nz.mem[390] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00365_) \MSYNC_1r1w.synth.nz.mem[391] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00366_) \MSYNC_1r1w.synth.nz.mem[392] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00367_) \MSYNC_1r1w.synth.nz.mem[393] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00368_) \MSYNC_1r1w.synth.nz.mem[394] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00369_) \MSYNC_1r1w.synth.nz.mem[395] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00370_) \MSYNC_1r1w.synth.nz.mem[396] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00371_) \MSYNC_1r1w.synth.nz.mem[397] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00372_) \MSYNC_1r1w.synth.nz.mem[398] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00375_) \MSYNC_1r1w.synth.nz.mem[3] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00376_) \MSYNC_1r1w.synth.nz.mem[400] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00377_) \MSYNC_1r1w.synth.nz.mem[401] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00378_) \MSYNC_1r1w.synth.nz.mem[402] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00379_) \MSYNC_1r1w.synth.nz.mem[403] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00380_) \MSYNC_1r1w.synth.nz.mem[404] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00381_) \MSYNC_1r1w.synth.nz.mem[405] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00382_) \MSYNC_1r1w.synth.nz.mem[406] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00383_) \MSYNC_1r1w.synth.nz.mem[407] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00384_) \MSYNC_1r1w.synth.nz.mem[408] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00386_) \MSYNC_1r1w.synth.nz.mem[40] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00387_) \MSYNC_1r1w.synth.nz.mem[410] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00388_) \MSYNC_1r1w.synth.nz.mem[411] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00389_) \MSYNC_1r1w.synth.nz.mem[412] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00390_) \MSYNC_1r1w.synth.nz.mem[413] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00391_) \MSYNC_1r1w.synth.nz.mem[414] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00392_) \MSYNC_1r1w.synth.nz.mem[415] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00393_) \MSYNC_1r1w.synth.nz.mem[416] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00394_) \MSYNC_1r1w.synth.nz.mem[417] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00395_) \MSYNC_1r1w.synth.nz.mem[418] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00397_) \MSYNC_1r1w.synth.nz.mem[41] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00398_) \MSYNC_1r1w.synth.nz.mem[420] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00399_) \MSYNC_1r1w.synth.nz.mem[421] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00400_) \MSYNC_1r1w.synth.nz.mem[422] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00401_) \MSYNC_1r1w.synth.nz.mem[423] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00402_) \MSYNC_1r1w.synth.nz.mem[424] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00403_) \MSYNC_1r1w.synth.nz.mem[425] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00404_) \MSYNC_1r1w.synth.nz.mem[426] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00405_) \MSYNC_1r1w.synth.nz.mem[427] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00406_) \MSYNC_1r1w.synth.nz.mem[428] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00408_) \MSYNC_1r1w.synth.nz.mem[42] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00409_) \MSYNC_1r1w.synth.nz.mem[430] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00410_) \MSYNC_1r1w.synth.nz.mem[431] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00411_) \MSYNC_1r1w.synth.nz.mem[432] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00412_) \MSYNC_1r1w.synth.nz.mem[433] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00413_) \MSYNC_1r1w.synth.nz.mem[434] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00414_) \MSYNC_1r1w.synth.nz.mem[435] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00415_) \MSYNC_1r1w.synth.nz.mem[436] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00416_) \MSYNC_1r1w.synth.nz.mem[437] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00417_) \MSYNC_1r1w.synth.nz.mem[438] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00419_) \MSYNC_1r1w.synth.nz.mem[43] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00420_) \MSYNC_1r1w.synth.nz.mem[440] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00421_) \MSYNC_1r1w.synth.nz.mem[441] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00422_) \MSYNC_1r1w.synth.nz.mem[442] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00423_) \MSYNC_1r1w.synth.nz.mem[443] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00424_) \MSYNC_1r1w.synth.nz.mem[444] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00425_) \MSYNC_1r1w.synth.nz.mem[445] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00426_) \MSYNC_1r1w.synth.nz.mem[446] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00427_) \MSYNC_1r1w.synth.nz.mem[447] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00428_) \MSYNC_1r1w.synth.nz.mem[448] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00430_) \MSYNC_1r1w.synth.nz.mem[44] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00431_) \MSYNC_1r1w.synth.nz.mem[450] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00432_) \MSYNC_1r1w.synth.nz.mem[451] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00433_) \MSYNC_1r1w.synth.nz.mem[452] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00434_) \MSYNC_1r1w.synth.nz.mem[453] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00435_) \MSYNC_1r1w.synth.nz.mem[454] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00436_) \MSYNC_1r1w.synth.nz.mem[455] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00437_) \MSYNC_1r1w.synth.nz.mem[456] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00438_) \MSYNC_1r1w.synth.nz.mem[457] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00439_) \MSYNC_1r1w.synth.nz.mem[458] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00441_) \MSYNC_1r1w.synth.nz.mem[45] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00442_) \MSYNC_1r1w.synth.nz.mem[460] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00443_) \MSYNC_1r1w.synth.nz.mem[461] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00444_) \MSYNC_1r1w.synth.nz.mem[462] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00445_) \MSYNC_1r1w.synth.nz.mem[463] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00446_) \MSYNC_1r1w.synth.nz.mem[464] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00447_) \MSYNC_1r1w.synth.nz.mem[465] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00448_) \MSYNC_1r1w.synth.nz.mem[466] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00449_) \MSYNC_1r1w.synth.nz.mem[467] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00450_) \MSYNC_1r1w.synth.nz.mem[468] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00452_) \MSYNC_1r1w.synth.nz.mem[46] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00453_) \MSYNC_1r1w.synth.nz.mem[470] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00454_) \MSYNC_1r1w.synth.nz.mem[471] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00455_) \MSYNC_1r1w.synth.nz.mem[472] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00456_) \MSYNC_1r1w.synth.nz.mem[473] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00457_) \MSYNC_1r1w.synth.nz.mem[474] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00458_) \MSYNC_1r1w.synth.nz.mem[475] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00459_) \MSYNC_1r1w.synth.nz.mem[476] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00460_) \MSYNC_1r1w.synth.nz.mem[477] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00461_) \MSYNC_1r1w.synth.nz.mem[478] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00463_) \MSYNC_1r1w.synth.nz.mem[47] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00464_) \MSYNC_1r1w.synth.nz.mem[480] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00465_) \MSYNC_1r1w.synth.nz.mem[481] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00466_) \MSYNC_1r1w.synth.nz.mem[482] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00467_) \MSYNC_1r1w.synth.nz.mem[483] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00468_) \MSYNC_1r1w.synth.nz.mem[484] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00469_) \MSYNC_1r1w.synth.nz.mem[485] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00470_) \MSYNC_1r1w.synth.nz.mem[486] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00471_) \MSYNC_1r1w.synth.nz.mem[487] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00472_) \MSYNC_1r1w.synth.nz.mem[488] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00474_) \MSYNC_1r1w.synth.nz.mem[48] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00475_) \MSYNC_1r1w.synth.nz.mem[490] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00476_) \MSYNC_1r1w.synth.nz.mem[491] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00477_) \MSYNC_1r1w.synth.nz.mem[492] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00478_) \MSYNC_1r1w.synth.nz.mem[493] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00479_) \MSYNC_1r1w.synth.nz.mem[494] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00480_) \MSYNC_1r1w.synth.nz.mem[495] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00481_) \MSYNC_1r1w.synth.nz.mem[496] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00482_) \MSYNC_1r1w.synth.nz.mem[497] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00483_) \MSYNC_1r1w.synth.nz.mem[498] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00486_) \MSYNC_1r1w.synth.nz.mem[4] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00487_) \MSYNC_1r1w.synth.nz.mem[500] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00488_) \MSYNC_1r1w.synth.nz.mem[501] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00489_) \MSYNC_1r1w.synth.nz.mem[502] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00490_) \MSYNC_1r1w.synth.nz.mem[503] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00491_) \MSYNC_1r1w.synth.nz.mem[504] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00492_) \MSYNC_1r1w.synth.nz.mem[505] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00493_) \MSYNC_1r1w.synth.nz.mem[506] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00494_) \MSYNC_1r1w.synth.nz.mem[507] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00495_) \MSYNC_1r1w.synth.nz.mem[508] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00497_) \MSYNC_1r1w.synth.nz.mem[50] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00498_) \MSYNC_1r1w.synth.nz.mem[510] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00499_) \MSYNC_1r1w.synth.nz.mem[511] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00500_) \MSYNC_1r1w.synth.nz.mem[512] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00501_) \MSYNC_1r1w.synth.nz.mem[513] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00502_) \MSYNC_1r1w.synth.nz.mem[514] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00503_) \MSYNC_1r1w.synth.nz.mem[515] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00504_) \MSYNC_1r1w.synth.nz.mem[516] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00505_) \MSYNC_1r1w.synth.nz.mem[517] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00506_) \MSYNC_1r1w.synth.nz.mem[518] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00508_) \MSYNC_1r1w.synth.nz.mem[51] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00509_) \MSYNC_1r1w.synth.nz.mem[520] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00510_) \MSYNC_1r1w.synth.nz.mem[521] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00511_) \MSYNC_1r1w.synth.nz.mem[522] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00512_) \MSYNC_1r1w.synth.nz.mem[523] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00513_) \MSYNC_1r1w.synth.nz.mem[524] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00514_) \MSYNC_1r1w.synth.nz.mem[525] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00515_) \MSYNC_1r1w.synth.nz.mem[526] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00516_) \MSYNC_1r1w.synth.nz.mem[527] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00517_) \MSYNC_1r1w.synth.nz.mem[528] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00519_) \MSYNC_1r1w.synth.nz.mem[52] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00520_) \MSYNC_1r1w.synth.nz.mem[530] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00521_) \MSYNC_1r1w.synth.nz.mem[531] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00522_) \MSYNC_1r1w.synth.nz.mem[532] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00523_) \MSYNC_1r1w.synth.nz.mem[533] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00524_) \MSYNC_1r1w.synth.nz.mem[534] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00525_) \MSYNC_1r1w.synth.nz.mem[535] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00526_) \MSYNC_1r1w.synth.nz.mem[536] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00527_) \MSYNC_1r1w.synth.nz.mem[537] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00528_) \MSYNC_1r1w.synth.nz.mem[538] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00530_) \MSYNC_1r1w.synth.nz.mem[53] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00531_) \MSYNC_1r1w.synth.nz.mem[540] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00532_) \MSYNC_1r1w.synth.nz.mem[541] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00533_) \MSYNC_1r1w.synth.nz.mem[542] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00534_) \MSYNC_1r1w.synth.nz.mem[543] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00535_) \MSYNC_1r1w.synth.nz.mem[544] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00536_) \MSYNC_1r1w.synth.nz.mem[545] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00537_) \MSYNC_1r1w.synth.nz.mem[546] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00538_) \MSYNC_1r1w.synth.nz.mem[547] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00539_) \MSYNC_1r1w.synth.nz.mem[548] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00541_) \MSYNC_1r1w.synth.nz.mem[54] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00542_) \MSYNC_1r1w.synth.nz.mem[550] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00543_) \MSYNC_1r1w.synth.nz.mem[551] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00544_) \MSYNC_1r1w.synth.nz.mem[552] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00545_) \MSYNC_1r1w.synth.nz.mem[553] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00546_) \MSYNC_1r1w.synth.nz.mem[554] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00547_) \MSYNC_1r1w.synth.nz.mem[555] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00548_) \MSYNC_1r1w.synth.nz.mem[556] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00549_) \MSYNC_1r1w.synth.nz.mem[557] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00550_) \MSYNC_1r1w.synth.nz.mem[558] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00552_) \MSYNC_1r1w.synth.nz.mem[55] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00553_) \MSYNC_1r1w.synth.nz.mem[560] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00554_) \MSYNC_1r1w.synth.nz.mem[561] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00555_) \MSYNC_1r1w.synth.nz.mem[562] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00556_) \MSYNC_1r1w.synth.nz.mem[563] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00557_) \MSYNC_1r1w.synth.nz.mem[564] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00558_) \MSYNC_1r1w.synth.nz.mem[565] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00559_) \MSYNC_1r1w.synth.nz.mem[566] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00560_) \MSYNC_1r1w.synth.nz.mem[567] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00561_) \MSYNC_1r1w.synth.nz.mem[568] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00563_) \MSYNC_1r1w.synth.nz.mem[56] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00564_) \MSYNC_1r1w.synth.nz.mem[570] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00565_) \MSYNC_1r1w.synth.nz.mem[571] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00566_) \MSYNC_1r1w.synth.nz.mem[572] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00567_) \MSYNC_1r1w.synth.nz.mem[573] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00568_) \MSYNC_1r1w.synth.nz.mem[574] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00569_) \MSYNC_1r1w.synth.nz.mem[575] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00570_) \MSYNC_1r1w.synth.nz.mem[576] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00571_) \MSYNC_1r1w.synth.nz.mem[577] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00572_) \MSYNC_1r1w.synth.nz.mem[578] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00574_) \MSYNC_1r1w.synth.nz.mem[57] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00575_) \MSYNC_1r1w.synth.nz.mem[580] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00576_) \MSYNC_1r1w.synth.nz.mem[581] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00577_) \MSYNC_1r1w.synth.nz.mem[582] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00578_) \MSYNC_1r1w.synth.nz.mem[583] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00579_) \MSYNC_1r1w.synth.nz.mem[584] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00580_) \MSYNC_1r1w.synth.nz.mem[585] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00581_) \MSYNC_1r1w.synth.nz.mem[586] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00582_) \MSYNC_1r1w.synth.nz.mem[587] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00583_) \MSYNC_1r1w.synth.nz.mem[588] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00585_) \MSYNC_1r1w.synth.nz.mem[58] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00586_) \MSYNC_1r1w.synth.nz.mem[590] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00587_) \MSYNC_1r1w.synth.nz.mem[591] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00588_) \MSYNC_1r1w.synth.nz.mem[592] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00589_) \MSYNC_1r1w.synth.nz.mem[593] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00590_) \MSYNC_1r1w.synth.nz.mem[594] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00591_) \MSYNC_1r1w.synth.nz.mem[595] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00592_) \MSYNC_1r1w.synth.nz.mem[596] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00593_) \MSYNC_1r1w.synth.nz.mem[597] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00594_) \MSYNC_1r1w.synth.nz.mem[598] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00597_) \MSYNC_1r1w.synth.nz.mem[5] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00598_) \MSYNC_1r1w.synth.nz.mem[600] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00599_) \MSYNC_1r1w.synth.nz.mem[601] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00600_) \MSYNC_1r1w.synth.nz.mem[602] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00601_) \MSYNC_1r1w.synth.nz.mem[603] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00602_) \MSYNC_1r1w.synth.nz.mem[604] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00603_) \MSYNC_1r1w.synth.nz.mem[605] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00604_) \MSYNC_1r1w.synth.nz.mem[606] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00605_) \MSYNC_1r1w.synth.nz.mem[607] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00606_) \MSYNC_1r1w.synth.nz.mem[608] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00608_) \MSYNC_1r1w.synth.nz.mem[60] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00609_) \MSYNC_1r1w.synth.nz.mem[610] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00610_) \MSYNC_1r1w.synth.nz.mem[611] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00611_) \MSYNC_1r1w.synth.nz.mem[612] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00612_) \MSYNC_1r1w.synth.nz.mem[613] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00613_) \MSYNC_1r1w.synth.nz.mem[614] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00614_) \MSYNC_1r1w.synth.nz.mem[615] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00615_) \MSYNC_1r1w.synth.nz.mem[616] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00616_) \MSYNC_1r1w.synth.nz.mem[617] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00617_) \MSYNC_1r1w.synth.nz.mem[618] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00619_) \MSYNC_1r1w.synth.nz.mem[61] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00620_) \MSYNC_1r1w.synth.nz.mem[620] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00621_) \MSYNC_1r1w.synth.nz.mem[621] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00622_) \MSYNC_1r1w.synth.nz.mem[622] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00623_) \MSYNC_1r1w.synth.nz.mem[623] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00624_) \MSYNC_1r1w.synth.nz.mem[624] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00625_) \MSYNC_1r1w.synth.nz.mem[625] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00626_) \MSYNC_1r1w.synth.nz.mem[626] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00627_) \MSYNC_1r1w.synth.nz.mem[627] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00628_) \MSYNC_1r1w.synth.nz.mem[628] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00630_) \MSYNC_1r1w.synth.nz.mem[62] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00631_) \MSYNC_1r1w.synth.nz.mem[630] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00632_) \MSYNC_1r1w.synth.nz.mem[631] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00633_) \MSYNC_1r1w.synth.nz.mem[632] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00634_) \MSYNC_1r1w.synth.nz.mem[633] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00635_) \MSYNC_1r1w.synth.nz.mem[634] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00636_) \MSYNC_1r1w.synth.nz.mem[635] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00637_) \MSYNC_1r1w.synth.nz.mem[636] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00638_) \MSYNC_1r1w.synth.nz.mem[637] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00639_) \MSYNC_1r1w.synth.nz.mem[638] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00641_) \MSYNC_1r1w.synth.nz.mem[63] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00642_) \MSYNC_1r1w.synth.nz.mem[640] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00643_) \MSYNC_1r1w.synth.nz.mem[641] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00644_) \MSYNC_1r1w.synth.nz.mem[642] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00645_) \MSYNC_1r1w.synth.nz.mem[643] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00646_) \MSYNC_1r1w.synth.nz.mem[644] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00647_) \MSYNC_1r1w.synth.nz.mem[645] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00648_) \MSYNC_1r1w.synth.nz.mem[646] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00649_) \MSYNC_1r1w.synth.nz.mem[647] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00650_) \MSYNC_1r1w.synth.nz.mem[648] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00652_) \MSYNC_1r1w.synth.nz.mem[64] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00653_) \MSYNC_1r1w.synth.nz.mem[650] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00654_) \MSYNC_1r1w.synth.nz.mem[651] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00655_) \MSYNC_1r1w.synth.nz.mem[652] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00656_) \MSYNC_1r1w.synth.nz.mem[653] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00657_) \MSYNC_1r1w.synth.nz.mem[654] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00658_) \MSYNC_1r1w.synth.nz.mem[655] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00659_) \MSYNC_1r1w.synth.nz.mem[656] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00660_) \MSYNC_1r1w.synth.nz.mem[657] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00661_) \MSYNC_1r1w.synth.nz.mem[658] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00663_) \MSYNC_1r1w.synth.nz.mem[65] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00664_) \MSYNC_1r1w.synth.nz.mem[660] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00665_) \MSYNC_1r1w.synth.nz.mem[661] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00666_) \MSYNC_1r1w.synth.nz.mem[662] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00667_) \MSYNC_1r1w.synth.nz.mem[663] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00668_) \MSYNC_1r1w.synth.nz.mem[664] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00669_) \MSYNC_1r1w.synth.nz.mem[665] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00670_) \MSYNC_1r1w.synth.nz.mem[666] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00671_) \MSYNC_1r1w.synth.nz.mem[667] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00672_) \MSYNC_1r1w.synth.nz.mem[668] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00674_) \MSYNC_1r1w.synth.nz.mem[66] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00675_) \MSYNC_1r1w.synth.nz.mem[670] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00676_) \MSYNC_1r1w.synth.nz.mem[671] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00677_) \MSYNC_1r1w.synth.nz.mem[672] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00678_) \MSYNC_1r1w.synth.nz.mem[673] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00679_) \MSYNC_1r1w.synth.nz.mem[674] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00680_) \MSYNC_1r1w.synth.nz.mem[675] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00681_) \MSYNC_1r1w.synth.nz.mem[676] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00682_) \MSYNC_1r1w.synth.nz.mem[677] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00683_) \MSYNC_1r1w.synth.nz.mem[678] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00685_) \MSYNC_1r1w.synth.nz.mem[67] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00686_) \MSYNC_1r1w.synth.nz.mem[680] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00687_) \MSYNC_1r1w.synth.nz.mem[681] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00688_) \MSYNC_1r1w.synth.nz.mem[682] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00689_) \MSYNC_1r1w.synth.nz.mem[683] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00690_) \MSYNC_1r1w.synth.nz.mem[684] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00691_) \MSYNC_1r1w.synth.nz.mem[685] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00692_) \MSYNC_1r1w.synth.nz.mem[686] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00693_) \MSYNC_1r1w.synth.nz.mem[687] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00694_) \MSYNC_1r1w.synth.nz.mem[688] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00696_) \MSYNC_1r1w.synth.nz.mem[68] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00697_) \MSYNC_1r1w.synth.nz.mem[690] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00698_) \MSYNC_1r1w.synth.nz.mem[691] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00699_) \MSYNC_1r1w.synth.nz.mem[692] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00700_) \MSYNC_1r1w.synth.nz.mem[693] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00701_) \MSYNC_1r1w.synth.nz.mem[694] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00702_) \MSYNC_1r1w.synth.nz.mem[695] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00703_) \MSYNC_1r1w.synth.nz.mem[696] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00704_) \MSYNC_1r1w.synth.nz.mem[697] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00705_) \MSYNC_1r1w.synth.nz.mem[698] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00708_) \MSYNC_1r1w.synth.nz.mem[6] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00709_) \MSYNC_1r1w.synth.nz.mem[700] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00710_) \MSYNC_1r1w.synth.nz.mem[701] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00711_) \MSYNC_1r1w.synth.nz.mem[702] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00712_) \MSYNC_1r1w.synth.nz.mem[703] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00713_) \MSYNC_1r1w.synth.nz.mem[704] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00714_) \MSYNC_1r1w.synth.nz.mem[705] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00715_) \MSYNC_1r1w.synth.nz.mem[706] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00716_) \MSYNC_1r1w.synth.nz.mem[707] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00717_) \MSYNC_1r1w.synth.nz.mem[708] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00719_) \MSYNC_1r1w.synth.nz.mem[70] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00720_) \MSYNC_1r1w.synth.nz.mem[710] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00721_) \MSYNC_1r1w.synth.nz.mem[711] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00722_) \MSYNC_1r1w.synth.nz.mem[712] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00723_) \MSYNC_1r1w.synth.nz.mem[713] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00724_) \MSYNC_1r1w.synth.nz.mem[714] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00725_) \MSYNC_1r1w.synth.nz.mem[715] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00726_) \MSYNC_1r1w.synth.nz.mem[716] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00727_) \MSYNC_1r1w.synth.nz.mem[717] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00728_) \MSYNC_1r1w.synth.nz.mem[718] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00730_) \MSYNC_1r1w.synth.nz.mem[71] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00731_) \MSYNC_1r1w.synth.nz.mem[720] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00732_) \MSYNC_1r1w.synth.nz.mem[721] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00733_) \MSYNC_1r1w.synth.nz.mem[722] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00734_) \MSYNC_1r1w.synth.nz.mem[723] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00735_) \MSYNC_1r1w.synth.nz.mem[724] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00736_) \MSYNC_1r1w.synth.nz.mem[725] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00737_) \MSYNC_1r1w.synth.nz.mem[726] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00738_) \MSYNC_1r1w.synth.nz.mem[727] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00739_) \MSYNC_1r1w.synth.nz.mem[728] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00741_) \MSYNC_1r1w.synth.nz.mem[72] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00742_) \MSYNC_1r1w.synth.nz.mem[730] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00743_) \MSYNC_1r1w.synth.nz.mem[731] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00744_) \MSYNC_1r1w.synth.nz.mem[732] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00745_) \MSYNC_1r1w.synth.nz.mem[733] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00746_) \MSYNC_1r1w.synth.nz.mem[734] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00747_) \MSYNC_1r1w.synth.nz.mem[735] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00748_) \MSYNC_1r1w.synth.nz.mem[736] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00749_) \MSYNC_1r1w.synth.nz.mem[737] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00750_) \MSYNC_1r1w.synth.nz.mem[738] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00752_) \MSYNC_1r1w.synth.nz.mem[73] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00753_) \MSYNC_1r1w.synth.nz.mem[740] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00754_) \MSYNC_1r1w.synth.nz.mem[741] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00755_) \MSYNC_1r1w.synth.nz.mem[742] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00756_) \MSYNC_1r1w.synth.nz.mem[743] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00757_) \MSYNC_1r1w.synth.nz.mem[744] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00758_) \MSYNC_1r1w.synth.nz.mem[745] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00759_) \MSYNC_1r1w.synth.nz.mem[746] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00760_) \MSYNC_1r1w.synth.nz.mem[747] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00761_) \MSYNC_1r1w.synth.nz.mem[748] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00763_) \MSYNC_1r1w.synth.nz.mem[74] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00764_) \MSYNC_1r1w.synth.nz.mem[750] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00765_) \MSYNC_1r1w.synth.nz.mem[751] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00766_) \MSYNC_1r1w.synth.nz.mem[752] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00767_) \MSYNC_1r1w.synth.nz.mem[753] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00768_) \MSYNC_1r1w.synth.nz.mem[754] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00769_) \MSYNC_1r1w.synth.nz.mem[755] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00770_) \MSYNC_1r1w.synth.nz.mem[756] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00771_) \MSYNC_1r1w.synth.nz.mem[757] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00772_) \MSYNC_1r1w.synth.nz.mem[758] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00774_) \MSYNC_1r1w.synth.nz.mem[75] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00775_) \MSYNC_1r1w.synth.nz.mem[760] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00776_) \MSYNC_1r1w.synth.nz.mem[761] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00777_) \MSYNC_1r1w.synth.nz.mem[762] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00778_) \MSYNC_1r1w.synth.nz.mem[763] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00779_) \MSYNC_1r1w.synth.nz.mem[764] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00780_) \MSYNC_1r1w.synth.nz.mem[765] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00781_) \MSYNC_1r1w.synth.nz.mem[766] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00782_) \MSYNC_1r1w.synth.nz.mem[767] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00783_) \MSYNC_1r1w.synth.nz.mem[768] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00785_) \MSYNC_1r1w.synth.nz.mem[76] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00786_) \MSYNC_1r1w.synth.nz.mem[770] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00787_) \MSYNC_1r1w.synth.nz.mem[771] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00788_) \MSYNC_1r1w.synth.nz.mem[772] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00789_) \MSYNC_1r1w.synth.nz.mem[773] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00790_) \MSYNC_1r1w.synth.nz.mem[774] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00791_) \MSYNC_1r1w.synth.nz.mem[775] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00792_) \MSYNC_1r1w.synth.nz.mem[776] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00793_) \MSYNC_1r1w.synth.nz.mem[777] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00794_) \MSYNC_1r1w.synth.nz.mem[778] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00796_) \MSYNC_1r1w.synth.nz.mem[77] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00797_) \MSYNC_1r1w.synth.nz.mem[780] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00798_) \MSYNC_1r1w.synth.nz.mem[781] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00799_) \MSYNC_1r1w.synth.nz.mem[782] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00800_) \MSYNC_1r1w.synth.nz.mem[783] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00801_) \MSYNC_1r1w.synth.nz.mem[784] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00802_) \MSYNC_1r1w.synth.nz.mem[785] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00803_) \MSYNC_1r1w.synth.nz.mem[786] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00804_) \MSYNC_1r1w.synth.nz.mem[787] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00805_) \MSYNC_1r1w.synth.nz.mem[788] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00807_) \MSYNC_1r1w.synth.nz.mem[78] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00808_) \MSYNC_1r1w.synth.nz.mem[790] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00809_) \MSYNC_1r1w.synth.nz.mem[791] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00810_) \MSYNC_1r1w.synth.nz.mem[792] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00811_) \MSYNC_1r1w.synth.nz.mem[793] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00812_) \MSYNC_1r1w.synth.nz.mem[794] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00813_) \MSYNC_1r1w.synth.nz.mem[795] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00814_) \MSYNC_1r1w.synth.nz.mem[796] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00815_) \MSYNC_1r1w.synth.nz.mem[797] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00816_) \MSYNC_1r1w.synth.nz.mem[798] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00819_) \MSYNC_1r1w.synth.nz.mem[7] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00820_) \MSYNC_1r1w.synth.nz.mem[800] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00821_) \MSYNC_1r1w.synth.nz.mem[801] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00822_) \MSYNC_1r1w.synth.nz.mem[802] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00823_) \MSYNC_1r1w.synth.nz.mem[803] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00824_) \MSYNC_1r1w.synth.nz.mem[804] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00825_) \MSYNC_1r1w.synth.nz.mem[805] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00826_) \MSYNC_1r1w.synth.nz.mem[806] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00827_) \MSYNC_1r1w.synth.nz.mem[807] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00828_) \MSYNC_1r1w.synth.nz.mem[808] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00830_) \MSYNC_1r1w.synth.nz.mem[80] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00831_) \MSYNC_1r1w.synth.nz.mem[810] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00832_) \MSYNC_1r1w.synth.nz.mem[811] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00833_) \MSYNC_1r1w.synth.nz.mem[812] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00834_) \MSYNC_1r1w.synth.nz.mem[813] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00835_) \MSYNC_1r1w.synth.nz.mem[814] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00836_) \MSYNC_1r1w.synth.nz.mem[815] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00837_) \MSYNC_1r1w.synth.nz.mem[816] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00838_) \MSYNC_1r1w.synth.nz.mem[817] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00839_) \MSYNC_1r1w.synth.nz.mem[818] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00841_) \MSYNC_1r1w.synth.nz.mem[81] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00842_) \MSYNC_1r1w.synth.nz.mem[820] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00843_) \MSYNC_1r1w.synth.nz.mem[821] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00844_) \MSYNC_1r1w.synth.nz.mem[822] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00845_) \MSYNC_1r1w.synth.nz.mem[823] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00846_) \MSYNC_1r1w.synth.nz.mem[824] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00847_) \MSYNC_1r1w.synth.nz.mem[825] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00848_) \MSYNC_1r1w.synth.nz.mem[826] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00849_) \MSYNC_1r1w.synth.nz.mem[827] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00850_) \MSYNC_1r1w.synth.nz.mem[828] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00852_) \MSYNC_1r1w.synth.nz.mem[82] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00853_) \MSYNC_1r1w.synth.nz.mem[830] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00854_) \MSYNC_1r1w.synth.nz.mem[831] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00855_) \MSYNC_1r1w.synth.nz.mem[832] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00856_) \MSYNC_1r1w.synth.nz.mem[833] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00857_) \MSYNC_1r1w.synth.nz.mem[834] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00858_) \MSYNC_1r1w.synth.nz.mem[835] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00859_) \MSYNC_1r1w.synth.nz.mem[836] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00860_) \MSYNC_1r1w.synth.nz.mem[837] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00861_) \MSYNC_1r1w.synth.nz.mem[838] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00863_) \MSYNC_1r1w.synth.nz.mem[83] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00864_) \MSYNC_1r1w.synth.nz.mem[840] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00865_) \MSYNC_1r1w.synth.nz.mem[841] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00866_) \MSYNC_1r1w.synth.nz.mem[842] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00867_) \MSYNC_1r1w.synth.nz.mem[843] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00868_) \MSYNC_1r1w.synth.nz.mem[844] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00869_) \MSYNC_1r1w.synth.nz.mem[845] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00870_) \MSYNC_1r1w.synth.nz.mem[846] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00871_) \MSYNC_1r1w.synth.nz.mem[847] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00872_) \MSYNC_1r1w.synth.nz.mem[848] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00874_) \MSYNC_1r1w.synth.nz.mem[84] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00875_) \MSYNC_1r1w.synth.nz.mem[850] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00876_) \MSYNC_1r1w.synth.nz.mem[851] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00877_) \MSYNC_1r1w.synth.nz.mem[852] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00878_) \MSYNC_1r1w.synth.nz.mem[853] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00879_) \MSYNC_1r1w.synth.nz.mem[854] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00880_) \MSYNC_1r1w.synth.nz.mem[855] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00881_) \MSYNC_1r1w.synth.nz.mem[856] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00882_) \MSYNC_1r1w.synth.nz.mem[857] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00883_) \MSYNC_1r1w.synth.nz.mem[858] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00885_) \MSYNC_1r1w.synth.nz.mem[85] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00886_) \MSYNC_1r1w.synth.nz.mem[860] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00887_) \MSYNC_1r1w.synth.nz.mem[861] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00888_) \MSYNC_1r1w.synth.nz.mem[862] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00889_) \MSYNC_1r1w.synth.nz.mem[863] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00890_) \MSYNC_1r1w.synth.nz.mem[864] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00891_) \MSYNC_1r1w.synth.nz.mem[865] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00892_) \MSYNC_1r1w.synth.nz.mem[866] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00893_) \MSYNC_1r1w.synth.nz.mem[867] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00894_) \MSYNC_1r1w.synth.nz.mem[868] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00896_) \MSYNC_1r1w.synth.nz.mem[86] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00897_) \MSYNC_1r1w.synth.nz.mem[870] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00898_) \MSYNC_1r1w.synth.nz.mem[871] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00899_) \MSYNC_1r1w.synth.nz.mem[872] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00900_) \MSYNC_1r1w.synth.nz.mem[873] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00901_) \MSYNC_1r1w.synth.nz.mem[874] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00902_) \MSYNC_1r1w.synth.nz.mem[875] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00903_) \MSYNC_1r1w.synth.nz.mem[876] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00904_) \MSYNC_1r1w.synth.nz.mem[877] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00905_) \MSYNC_1r1w.synth.nz.mem[878] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00907_) \MSYNC_1r1w.synth.nz.mem[87] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00908_) \MSYNC_1r1w.synth.nz.mem[880] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00909_) \MSYNC_1r1w.synth.nz.mem[881] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00910_) \MSYNC_1r1w.synth.nz.mem[882] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00911_) \MSYNC_1r1w.synth.nz.mem[883] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00912_) \MSYNC_1r1w.synth.nz.mem[884] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00913_) \MSYNC_1r1w.synth.nz.mem[885] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00914_) \MSYNC_1r1w.synth.nz.mem[886] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00915_) \MSYNC_1r1w.synth.nz.mem[887] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00916_) \MSYNC_1r1w.synth.nz.mem[888] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00918_) \MSYNC_1r1w.synth.nz.mem[88] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00919_) \MSYNC_1r1w.synth.nz.mem[890] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00920_) \MSYNC_1r1w.synth.nz.mem[891] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00921_) \MSYNC_1r1w.synth.nz.mem[892] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00922_) \MSYNC_1r1w.synth.nz.mem[893] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00923_) \MSYNC_1r1w.synth.nz.mem[894] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00924_) \MSYNC_1r1w.synth.nz.mem[895] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00925_) \MSYNC_1r1w.synth.nz.mem[896] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00926_) \MSYNC_1r1w.synth.nz.mem[897] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00927_) \MSYNC_1r1w.synth.nz.mem[898] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00930_) \MSYNC_1r1w.synth.nz.mem[8] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00931_) \MSYNC_1r1w.synth.nz.mem[900] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00932_) \MSYNC_1r1w.synth.nz.mem[901] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00933_) \MSYNC_1r1w.synth.nz.mem[902] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00934_) \MSYNC_1r1w.synth.nz.mem[903] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00935_) \MSYNC_1r1w.synth.nz.mem[904] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00936_) \MSYNC_1r1w.synth.nz.mem[905] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00937_) \MSYNC_1r1w.synth.nz.mem[906] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00938_) \MSYNC_1r1w.synth.nz.mem[907] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00939_) \MSYNC_1r1w.synth.nz.mem[908] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00941_) \MSYNC_1r1w.synth.nz.mem[90] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00942_) \MSYNC_1r1w.synth.nz.mem[910] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00943_) \MSYNC_1r1w.synth.nz.mem[911] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00944_) \MSYNC_1r1w.synth.nz.mem[912] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00945_) \MSYNC_1r1w.synth.nz.mem[913] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00946_) \MSYNC_1r1w.synth.nz.mem[914] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00947_) \MSYNC_1r1w.synth.nz.mem[915] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00948_) \MSYNC_1r1w.synth.nz.mem[916] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00949_) \MSYNC_1r1w.synth.nz.mem[917] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00950_) \MSYNC_1r1w.synth.nz.mem[918] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00952_) \MSYNC_1r1w.synth.nz.mem[91] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00953_) \MSYNC_1r1w.synth.nz.mem[920] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00954_) \MSYNC_1r1w.synth.nz.mem[921] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00955_) \MSYNC_1r1w.synth.nz.mem[922] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00956_) \MSYNC_1r1w.synth.nz.mem[923] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00957_) \MSYNC_1r1w.synth.nz.mem[924] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00958_) \MSYNC_1r1w.synth.nz.mem[925] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00959_) \MSYNC_1r1w.synth.nz.mem[926] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00960_) \MSYNC_1r1w.synth.nz.mem[927] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00961_) \MSYNC_1r1w.synth.nz.mem[928] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00963_) \MSYNC_1r1w.synth.nz.mem[92] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00964_) \MSYNC_1r1w.synth.nz.mem[930] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00965_) \MSYNC_1r1w.synth.nz.mem[931] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00966_) \MSYNC_1r1w.synth.nz.mem[932] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00967_) \MSYNC_1r1w.synth.nz.mem[933] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00968_) \MSYNC_1r1w.synth.nz.mem[934] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00969_) \MSYNC_1r1w.synth.nz.mem[935] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00970_) \MSYNC_1r1w.synth.nz.mem[936] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00971_) \MSYNC_1r1w.synth.nz.mem[937] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00972_) \MSYNC_1r1w.synth.nz.mem[938] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00974_) \MSYNC_1r1w.synth.nz.mem[93] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00975_) \MSYNC_1r1w.synth.nz.mem[940] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00976_) \MSYNC_1r1w.synth.nz.mem[941] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00977_) \MSYNC_1r1w.synth.nz.mem[942] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00978_) \MSYNC_1r1w.synth.nz.mem[943] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00979_) \MSYNC_1r1w.synth.nz.mem[944] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00980_) \MSYNC_1r1w.synth.nz.mem[945] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00981_) \MSYNC_1r1w.synth.nz.mem[946] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00982_) \MSYNC_1r1w.synth.nz.mem[947] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00983_) \MSYNC_1r1w.synth.nz.mem[948] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00985_) \MSYNC_1r1w.synth.nz.mem[94] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00986_) \MSYNC_1r1w.synth.nz.mem[950] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00987_) \MSYNC_1r1w.synth.nz.mem[951] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00988_) \MSYNC_1r1w.synth.nz.mem[952] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00989_) \MSYNC_1r1w.synth.nz.mem[953] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00990_) \MSYNC_1r1w.synth.nz.mem[954] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00991_) \MSYNC_1r1w.synth.nz.mem[955] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00992_) \MSYNC_1r1w.synth.nz.mem[956] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00993_) \MSYNC_1r1w.synth.nz.mem[957] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00994_) \MSYNC_1r1w.synth.nz.mem[958] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00996_) \MSYNC_1r1w.synth.nz.mem[95] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00997_) \MSYNC_1r1w.synth.nz.mem[960] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00998_) \MSYNC_1r1w.synth.nz.mem[961] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00999_) \MSYNC_1r1w.synth.nz.mem[962] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01000_) \MSYNC_1r1w.synth.nz.mem[963] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01001_) \MSYNC_1r1w.synth.nz.mem[964] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01002_) \MSYNC_1r1w.synth.nz.mem[965] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01003_) \MSYNC_1r1w.synth.nz.mem[966] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01004_) \MSYNC_1r1w.synth.nz.mem[967] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01005_) \MSYNC_1r1w.synth.nz.mem[968] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01007_) \MSYNC_1r1w.synth.nz.mem[96] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01008_) \MSYNC_1r1w.synth.nz.mem[970] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01009_) \MSYNC_1r1w.synth.nz.mem[971] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01010_) \MSYNC_1r1w.synth.nz.mem[972] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01011_) \MSYNC_1r1w.synth.nz.mem[973] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01012_) \MSYNC_1r1w.synth.nz.mem[974] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01013_) \MSYNC_1r1w.synth.nz.mem[975] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01014_) \MSYNC_1r1w.synth.nz.mem[976] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01015_) \MSYNC_1r1w.synth.nz.mem[977] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01016_) \MSYNC_1r1w.synth.nz.mem[978] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01018_) \MSYNC_1r1w.synth.nz.mem[97] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01019_) \MSYNC_1r1w.synth.nz.mem[980] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01020_) \MSYNC_1r1w.synth.nz.mem[981] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01021_) \MSYNC_1r1w.synth.nz.mem[982] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01022_) \MSYNC_1r1w.synth.nz.mem[983] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01023_) \MSYNC_1r1w.synth.nz.mem[984] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01024_) \MSYNC_1r1w.synth.nz.mem[985] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01025_) \MSYNC_1r1w.synth.nz.mem[986] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01026_) \MSYNC_1r1w.synth.nz.mem[987] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01027_) \MSYNC_1r1w.synth.nz.mem[988] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01029_) \MSYNC_1r1w.synth.nz.mem[98] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01030_) \MSYNC_1r1w.synth.nz.mem[990] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01031_) \MSYNC_1r1w.synth.nz.mem[991] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01032_) \MSYNC_1r1w.synth.nz.mem[992] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01033_) \MSYNC_1r1w.synth.nz.mem[993] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01034_) \MSYNC_1r1w.synth.nz.mem[994] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01035_) \MSYNC_1r1w.synth.nz.mem[995] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01036_) \MSYNC_1r1w.synth.nz.mem[996] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01037_) \MSYNC_1r1w.synth.nz.mem[997] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01038_) \MSYNC_1r1w.synth.nz.mem[998] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00018_) \MSYNC_1r1w.synth.nz.mem[0] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00019_) \MSYNC_1r1w.synth.nz.mem[1000] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00020_) \MSYNC_1r1w.synth.nz.mem[1001] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00021_) \MSYNC_1r1w.synth.nz.mem[1002] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00022_) \MSYNC_1r1w.synth.nz.mem[1003] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00023_) \MSYNC_1r1w.synth.nz.mem[1004] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00024_) \MSYNC_1r1w.synth.nz.mem[1005] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00025_) \MSYNC_1r1w.synth.nz.mem[1006] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00026_) \MSYNC_1r1w.synth.nz.mem[1007] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00027_) \MSYNC_1r1w.synth.nz.mem[1008] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00029_) \MSYNC_1r1w.synth.nz.mem[100] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00030_) \MSYNC_1r1w.synth.nz.mem[1010] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00031_) \MSYNC_1r1w.synth.nz.mem[1011] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00032_) \MSYNC_1r1w.synth.nz.mem[1012] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00033_) \MSYNC_1r1w.synth.nz.mem[1013] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00034_) \MSYNC_1r1w.synth.nz.mem[1014] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00035_) \MSYNC_1r1w.synth.nz.mem[1015] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00036_) \MSYNC_1r1w.synth.nz.mem[1016] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00037_) \MSYNC_1r1w.synth.nz.mem[1017] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00038_) \MSYNC_1r1w.synth.nz.mem[1018] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00040_) \MSYNC_1r1w.synth.nz.mem[101] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00041_) \MSYNC_1r1w.synth.nz.mem[1020] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00042_) \MSYNC_1r1w.synth.nz.mem[1021] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_00043_) \MSYNC_1r1w.synth.nz.mem[1022] [15] <= w_data_i[15];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [0] <= w_data_i[0];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [1] <= w_data_i[1];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [2] <= w_data_i[2];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [3] <= w_data_i[3];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [4] <= w_data_i[4];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [5] <= w_data_i[5];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [6] <= w_data_i[6];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [7] <= w_data_i[7];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [8] <= w_data_i[8];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [9] <= w_data_i[9];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [10] <= w_data_i[10];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [11] <= w_data_i[11];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [12] <= w_data_i[12];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [13] <= w_data_i[13];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [14] <= w_data_i[14];
  always @(posedge w_clk_i)
    if (_01041_) \MSYNC_1r1w.synth.nz.mem[9] [15] <= w_data_i[15];
  assign \MSYNC_1r1w.r_addr_i  = \bapg_rd.w_ptr_r [9:0];
  assign \MSYNC_1r1w.r_data_o  = r_data_o;
  assign \MSYNC_1r1w.r_v_i  = r_valid_o;
  assign \MSYNC_1r1w.synth.r_addr_i  = \bapg_rd.w_ptr_r [9:0];
  assign \MSYNC_1r1w.synth.r_data_o  = r_data_o;
  assign \MSYNC_1r1w.synth.r_v_i  = r_valid_o;
  assign \MSYNC_1r1w.synth.unused0  = w_reset_i;
  assign \MSYNC_1r1w.synth.unused1  = r_valid_o;
  assign \MSYNC_1r1w.synth.w_addr_i  = \bapg_wr.w_ptr_r [9:0];
  assign \MSYNC_1r1w.synth.w_clk_i  = w_clk_i;
  assign \MSYNC_1r1w.synth.w_data_i  = w_data_i;
  assign \MSYNC_1r1w.synth.w_reset_i  = w_reset_i;
  assign \MSYNC_1r1w.synth.w_v_i  = w_enq_i;
  assign \MSYNC_1r1w.w_addr_i  = \bapg_wr.w_ptr_r [9:0];
  assign \MSYNC_1r1w.w_clk_i  = w_clk_i;
  assign \MSYNC_1r1w.w_data_i  = w_data_i;
  assign \MSYNC_1r1w.w_reset_i  = w_reset_i;
  assign \MSYNC_1r1w.w_v_i  = w_enq_i;
  assign \bapg_rd.ptr_sync.iclk_data_o  = { \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r , \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_rd.w_ptr_p1_r [1] };
  assign \bapg_rd.ptr_sync.iclk_i  = r_clk_i;
  assign \bapg_rd.ptr_sync.iclk_reset_i  = r_reset_i;
  assign \bapg_rd.ptr_sync.oclk_data_o  = { \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r , \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r  };
  assign \bapg_rd.ptr_sync.oclk_i  = w_clk_i;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [0] = \bapg_rd.w_ptr_p1_r [1];
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.iclk_data_o  = { \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_rd.w_ptr_p1_r [1] };
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.iclk_i  = r_clk_i;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.iclk_reset_i  = r_reset_i;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.oclk_data_o  = \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r ;
  assign \bapg_rd.ptr_sync.sync.p.maxb[0].blss.oclk_i  = w_clk_i;
  assign \bapg_rd.ptr_sync.sync.p.z.blss.iclk_data_o  = \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \bapg_rd.ptr_sync.sync.p.z.blss.iclk_i  = r_clk_i;
  assign \bapg_rd.ptr_sync.sync.p.z.blss.iclk_reset_i  = r_reset_i;
  assign \bapg_rd.ptr_sync.sync.p.z.blss.oclk_data_o  = \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \bapg_rd.ptr_sync.sync.p.z.blss.oclk_i  = w_clk_i;
  assign \bapg_rd.r_clk_i  = w_clk_i;
  assign \bapg_rd.w_clk_i  = r_clk_i;
  assign \bapg_rd.w_inc_i  = r_deq_i;
  assign \bapg_rd.w_ptr_binary_r_o  = { 1'hx, \bapg_rd.w_ptr_r [9:0] };
  assign \bapg_rd.w_ptr_gray_r  = { \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r , \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_rd.w_ptr_p1_r [1] };
  assign \bapg_rd.w_ptr_gray_r_o  = { \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r , \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_rd.w_ptr_p1_r [1] };
  assign \bapg_rd.w_ptr_gray_r_rsync  = { \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r , \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r  };
  assign \bapg_rd.w_ptr_gray_r_rsync_o  = { \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r , \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r  };
  assign \bapg_rd.w_ptr_r [10] = 1'hx;
  assign \bapg_rd.w_reset_i  = r_reset_i;
  assign \bapg_wr.ptr_sync.iclk_data_o  = { \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r , \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_wr.w_ptr_p1_r [1] };
  assign \bapg_wr.ptr_sync.iclk_i  = w_clk_i;
  assign \bapg_wr.ptr_sync.iclk_reset_i  = w_reset_i;
  assign \bapg_wr.ptr_sync.oclk_data_o  = { \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r , \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r  };
  assign \bapg_wr.ptr_sync.oclk_i  = r_clk_i;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [0] = \bapg_wr.w_ptr_p1_r [1];
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.iclk_data_o  = { \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_wr.w_ptr_p1_r [1] };
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.iclk_i  = w_clk_i;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.iclk_reset_i  = w_reset_i;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.oclk_data_o  = \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r ;
  assign \bapg_wr.ptr_sync.sync.p.maxb[0].blss.oclk_i  = r_clk_i;
  assign \bapg_wr.ptr_sync.sync.p.z.blss.iclk_data_o  = \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r ;
  assign \bapg_wr.ptr_sync.sync.p.z.blss.iclk_i  = w_clk_i;
  assign \bapg_wr.ptr_sync.sync.p.z.blss.iclk_reset_i  = w_reset_i;
  assign \bapg_wr.ptr_sync.sync.p.z.blss.oclk_data_o  = \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r ;
  assign \bapg_wr.ptr_sync.sync.p.z.blss.oclk_i  = r_clk_i;
  assign \bapg_wr.r_clk_i  = r_clk_i;
  assign \bapg_wr.w_clk_i  = w_clk_i;
  assign \bapg_wr.w_inc_i  = w_enq_i;
  assign \bapg_wr.w_ptr_binary_r_o  = { 1'hx, \bapg_wr.w_ptr_r [9:0] };
  assign \bapg_wr.w_ptr_gray_r  = { \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r , \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_wr.w_ptr_p1_r [1] };
  assign \bapg_wr.w_ptr_gray_r_o  = { \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r , \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_wr.w_ptr_p1_r [1] };
  assign \bapg_wr.w_ptr_gray_r_rsync  = { \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r , \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r  };
  assign \bapg_wr.w_ptr_gray_r_rsync_o  = { \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r , \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r  };
  assign \bapg_wr.w_ptr_r [10] = 1'hx;
  assign \bapg_wr.w_reset_i  = w_reset_i;
  assign r_data_o_tmp = r_data_o;
  assign r_ptr_binary_r = { 1'hx, \bapg_rd.w_ptr_r [9:0] };
  assign r_ptr_gray_r = { \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r , \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_rd.w_ptr_p1_r [1] };
  assign r_ptr_gray_r_wsync = { \bapg_rd.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r , \bapg_rd.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r  };
  assign r_valid_o_tmp = r_valid_o;
  assign w_ptr_binary_r = { 1'hx, \bapg_wr.w_ptr_r [9:0] };
  assign w_ptr_gray_r = { \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_LNCH_r , \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_LNCH_r [7:1], \bapg_wr.w_ptr_p1_r [1] };
  assign w_ptr_gray_r_rsync = { \bapg_wr.ptr_sync.sync.p.z.blss.bsg_SYNC_2_r , \bapg_wr.ptr_sync.sync.p.maxb[0].blss.bsg_SYNC_2_r  };
endmodule
